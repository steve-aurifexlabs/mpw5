magic
tech sky130A
magscale 1 2
timestamp 1647896588
<< obsli1 >>
rect 1104 2159 238832 237745
<< obsm1 >>
rect 658 8 239738 237924
<< metal2 >>
rect 1030 239200 1086 240000
rect 3054 239200 3110 240000
rect 5170 239200 5226 240000
rect 7286 239200 7342 240000
rect 9402 239200 9458 240000
rect 11518 239200 11574 240000
rect 13634 239200 13690 240000
rect 15750 239200 15806 240000
rect 17866 239200 17922 240000
rect 19890 239200 19946 240000
rect 22006 239200 22062 240000
rect 24122 239200 24178 240000
rect 26238 239200 26294 240000
rect 28354 239200 28410 240000
rect 30470 239200 30526 240000
rect 32586 239200 32642 240000
rect 34702 239200 34758 240000
rect 36818 239200 36874 240000
rect 38842 239200 38898 240000
rect 40958 239200 41014 240000
rect 43074 239200 43130 240000
rect 45190 239200 45246 240000
rect 47306 239200 47362 240000
rect 49422 239200 49478 240000
rect 51538 239200 51594 240000
rect 53654 239200 53710 240000
rect 55770 239200 55826 240000
rect 57794 239200 57850 240000
rect 59910 239200 59966 240000
rect 62026 239200 62082 240000
rect 64142 239200 64198 240000
rect 66258 239200 66314 240000
rect 68374 239200 68430 240000
rect 70490 239200 70546 240000
rect 72606 239200 72662 240000
rect 74722 239200 74778 240000
rect 76746 239200 76802 240000
rect 78862 239200 78918 240000
rect 80978 239200 81034 240000
rect 83094 239200 83150 240000
rect 85210 239200 85266 240000
rect 87326 239200 87382 240000
rect 89442 239200 89498 240000
rect 91558 239200 91614 240000
rect 93582 239200 93638 240000
rect 95698 239200 95754 240000
rect 97814 239200 97870 240000
rect 99930 239200 99986 240000
rect 102046 239200 102102 240000
rect 104162 239200 104218 240000
rect 106278 239200 106334 240000
rect 108394 239200 108450 240000
rect 110510 239200 110566 240000
rect 112534 239200 112590 240000
rect 114650 239200 114706 240000
rect 116766 239200 116822 240000
rect 118882 239200 118938 240000
rect 120998 239200 121054 240000
rect 123114 239200 123170 240000
rect 125230 239200 125286 240000
rect 127346 239200 127402 240000
rect 129462 239200 129518 240000
rect 131486 239200 131542 240000
rect 133602 239200 133658 240000
rect 135718 239200 135774 240000
rect 137834 239200 137890 240000
rect 139950 239200 140006 240000
rect 142066 239200 142122 240000
rect 144182 239200 144238 240000
rect 146298 239200 146354 240000
rect 148414 239200 148470 240000
rect 150438 239200 150494 240000
rect 152554 239200 152610 240000
rect 154670 239200 154726 240000
rect 156786 239200 156842 240000
rect 158902 239200 158958 240000
rect 161018 239200 161074 240000
rect 163134 239200 163190 240000
rect 165250 239200 165306 240000
rect 167274 239200 167330 240000
rect 169390 239200 169446 240000
rect 171506 239200 171562 240000
rect 173622 239200 173678 240000
rect 175738 239200 175794 240000
rect 177854 239200 177910 240000
rect 179970 239200 180026 240000
rect 182086 239200 182142 240000
rect 184202 239200 184258 240000
rect 186226 239200 186282 240000
rect 188342 239200 188398 240000
rect 190458 239200 190514 240000
rect 192574 239200 192630 240000
rect 194690 239200 194746 240000
rect 196806 239200 196862 240000
rect 198922 239200 198978 240000
rect 201038 239200 201094 240000
rect 203154 239200 203210 240000
rect 205178 239200 205234 240000
rect 207294 239200 207350 240000
rect 209410 239200 209466 240000
rect 211526 239200 211582 240000
rect 213642 239200 213698 240000
rect 215758 239200 215814 240000
rect 217874 239200 217930 240000
rect 219990 239200 220046 240000
rect 222106 239200 222162 240000
rect 224130 239200 224186 240000
rect 226246 239200 226302 240000
rect 228362 239200 228418 240000
rect 230478 239200 230534 240000
rect 232594 239200 232650 240000
rect 234710 239200 234766 240000
rect 236826 239200 236882 240000
rect 238942 239200 238998 240000
rect 202 0 258 800
rect 662 0 718 800
rect 1122 0 1178 800
rect 1582 0 1638 800
rect 2134 0 2190 800
rect 2594 0 2650 800
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4066 0 4122 800
rect 4526 0 4582 800
rect 4986 0 5042 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7470 0 7526 800
rect 7930 0 7986 800
rect 8390 0 8446 800
rect 8942 0 8998 800
rect 9402 0 9458 800
rect 9862 0 9918 800
rect 10414 0 10470 800
rect 10874 0 10930 800
rect 11334 0 11390 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12806 0 12862 800
rect 13266 0 13322 800
rect 13818 0 13874 800
rect 14278 0 14334 800
rect 14738 0 14794 800
rect 15290 0 15346 800
rect 15750 0 15806 800
rect 16210 0 16266 800
rect 16670 0 16726 800
rect 17222 0 17278 800
rect 17682 0 17738 800
rect 18142 0 18198 800
rect 18694 0 18750 800
rect 19154 0 19210 800
rect 19614 0 19670 800
rect 20074 0 20130 800
rect 20626 0 20682 800
rect 21086 0 21142 800
rect 21546 0 21602 800
rect 22098 0 22154 800
rect 22558 0 22614 800
rect 23018 0 23074 800
rect 23570 0 23626 800
rect 24030 0 24086 800
rect 24490 0 24546 800
rect 24950 0 25006 800
rect 25502 0 25558 800
rect 25962 0 26018 800
rect 26422 0 26478 800
rect 26974 0 27030 800
rect 27434 0 27490 800
rect 27894 0 27950 800
rect 28354 0 28410 800
rect 28906 0 28962 800
rect 29366 0 29422 800
rect 29826 0 29882 800
rect 30378 0 30434 800
rect 30838 0 30894 800
rect 31298 0 31354 800
rect 31758 0 31814 800
rect 32310 0 32366 800
rect 32770 0 32826 800
rect 33230 0 33286 800
rect 33782 0 33838 800
rect 34242 0 34298 800
rect 34702 0 34758 800
rect 35254 0 35310 800
rect 35714 0 35770 800
rect 36174 0 36230 800
rect 36634 0 36690 800
rect 37186 0 37242 800
rect 37646 0 37702 800
rect 38106 0 38162 800
rect 38658 0 38714 800
rect 39118 0 39174 800
rect 39578 0 39634 800
rect 40038 0 40094 800
rect 40590 0 40646 800
rect 41050 0 41106 800
rect 41510 0 41566 800
rect 42062 0 42118 800
rect 42522 0 42578 800
rect 42982 0 43038 800
rect 43442 0 43498 800
rect 43994 0 44050 800
rect 44454 0 44510 800
rect 44914 0 44970 800
rect 45466 0 45522 800
rect 45926 0 45982 800
rect 46386 0 46442 800
rect 46938 0 46994 800
rect 47398 0 47454 800
rect 47858 0 47914 800
rect 48318 0 48374 800
rect 48870 0 48926 800
rect 49330 0 49386 800
rect 49790 0 49846 800
rect 50342 0 50398 800
rect 50802 0 50858 800
rect 51262 0 51318 800
rect 51722 0 51778 800
rect 52274 0 52330 800
rect 52734 0 52790 800
rect 53194 0 53250 800
rect 53746 0 53802 800
rect 54206 0 54262 800
rect 54666 0 54722 800
rect 55218 0 55274 800
rect 55678 0 55734 800
rect 56138 0 56194 800
rect 56598 0 56654 800
rect 57150 0 57206 800
rect 57610 0 57666 800
rect 58070 0 58126 800
rect 58622 0 58678 800
rect 59082 0 59138 800
rect 59542 0 59598 800
rect 60002 0 60058 800
rect 60554 0 60610 800
rect 61014 0 61070 800
rect 61474 0 61530 800
rect 62026 0 62082 800
rect 62486 0 62542 800
rect 62946 0 63002 800
rect 63406 0 63462 800
rect 63958 0 64014 800
rect 64418 0 64474 800
rect 64878 0 64934 800
rect 65430 0 65486 800
rect 65890 0 65946 800
rect 66350 0 66406 800
rect 66902 0 66958 800
rect 67362 0 67418 800
rect 67822 0 67878 800
rect 68282 0 68338 800
rect 68834 0 68890 800
rect 69294 0 69350 800
rect 69754 0 69810 800
rect 70306 0 70362 800
rect 70766 0 70822 800
rect 71226 0 71282 800
rect 71686 0 71742 800
rect 72238 0 72294 800
rect 72698 0 72754 800
rect 73158 0 73214 800
rect 73710 0 73766 800
rect 74170 0 74226 800
rect 74630 0 74686 800
rect 75090 0 75146 800
rect 75642 0 75698 800
rect 76102 0 76158 800
rect 76562 0 76618 800
rect 77114 0 77170 800
rect 77574 0 77630 800
rect 78034 0 78090 800
rect 78586 0 78642 800
rect 79046 0 79102 800
rect 79506 0 79562 800
rect 79966 0 80022 800
rect 80518 0 80574 800
rect 80978 0 81034 800
rect 81438 0 81494 800
rect 81990 0 82046 800
rect 82450 0 82506 800
rect 82910 0 82966 800
rect 83370 0 83426 800
rect 83922 0 83978 800
rect 84382 0 84438 800
rect 84842 0 84898 800
rect 85394 0 85450 800
rect 85854 0 85910 800
rect 86314 0 86370 800
rect 86774 0 86830 800
rect 87326 0 87382 800
rect 87786 0 87842 800
rect 88246 0 88302 800
rect 88798 0 88854 800
rect 89258 0 89314 800
rect 89718 0 89774 800
rect 90270 0 90326 800
rect 90730 0 90786 800
rect 91190 0 91246 800
rect 91650 0 91706 800
rect 92202 0 92258 800
rect 92662 0 92718 800
rect 93122 0 93178 800
rect 93674 0 93730 800
rect 94134 0 94190 800
rect 94594 0 94650 800
rect 95054 0 95110 800
rect 95606 0 95662 800
rect 96066 0 96122 800
rect 96526 0 96582 800
rect 97078 0 97134 800
rect 97538 0 97594 800
rect 97998 0 98054 800
rect 98550 0 98606 800
rect 99010 0 99066 800
rect 99470 0 99526 800
rect 99930 0 99986 800
rect 100482 0 100538 800
rect 100942 0 100998 800
rect 101402 0 101458 800
rect 101954 0 102010 800
rect 102414 0 102470 800
rect 102874 0 102930 800
rect 103334 0 103390 800
rect 103886 0 103942 800
rect 104346 0 104402 800
rect 104806 0 104862 800
rect 105358 0 105414 800
rect 105818 0 105874 800
rect 106278 0 106334 800
rect 106738 0 106794 800
rect 107290 0 107346 800
rect 107750 0 107806 800
rect 108210 0 108266 800
rect 108762 0 108818 800
rect 109222 0 109278 800
rect 109682 0 109738 800
rect 110234 0 110290 800
rect 110694 0 110750 800
rect 111154 0 111210 800
rect 111614 0 111670 800
rect 112166 0 112222 800
rect 112626 0 112682 800
rect 113086 0 113142 800
rect 113638 0 113694 800
rect 114098 0 114154 800
rect 114558 0 114614 800
rect 115018 0 115074 800
rect 115570 0 115626 800
rect 116030 0 116086 800
rect 116490 0 116546 800
rect 117042 0 117098 800
rect 117502 0 117558 800
rect 117962 0 118018 800
rect 118422 0 118478 800
rect 118974 0 119030 800
rect 119434 0 119490 800
rect 119894 0 119950 800
rect 120446 0 120502 800
rect 120906 0 120962 800
rect 121366 0 121422 800
rect 121918 0 121974 800
rect 122378 0 122434 800
rect 122838 0 122894 800
rect 123298 0 123354 800
rect 123850 0 123906 800
rect 124310 0 124366 800
rect 124770 0 124826 800
rect 125322 0 125378 800
rect 125782 0 125838 800
rect 126242 0 126298 800
rect 126702 0 126758 800
rect 127254 0 127310 800
rect 127714 0 127770 800
rect 128174 0 128230 800
rect 128726 0 128782 800
rect 129186 0 129242 800
rect 129646 0 129702 800
rect 130106 0 130162 800
rect 130658 0 130714 800
rect 131118 0 131174 800
rect 131578 0 131634 800
rect 132130 0 132186 800
rect 132590 0 132646 800
rect 133050 0 133106 800
rect 133602 0 133658 800
rect 134062 0 134118 800
rect 134522 0 134578 800
rect 134982 0 135038 800
rect 135534 0 135590 800
rect 135994 0 136050 800
rect 136454 0 136510 800
rect 137006 0 137062 800
rect 137466 0 137522 800
rect 137926 0 137982 800
rect 138386 0 138442 800
rect 138938 0 138994 800
rect 139398 0 139454 800
rect 139858 0 139914 800
rect 140410 0 140466 800
rect 140870 0 140926 800
rect 141330 0 141386 800
rect 141790 0 141846 800
rect 142342 0 142398 800
rect 142802 0 142858 800
rect 143262 0 143318 800
rect 143814 0 143870 800
rect 144274 0 144330 800
rect 144734 0 144790 800
rect 145286 0 145342 800
rect 145746 0 145802 800
rect 146206 0 146262 800
rect 146666 0 146722 800
rect 147218 0 147274 800
rect 147678 0 147734 800
rect 148138 0 148194 800
rect 148690 0 148746 800
rect 149150 0 149206 800
rect 149610 0 149666 800
rect 150070 0 150126 800
rect 150622 0 150678 800
rect 151082 0 151138 800
rect 151542 0 151598 800
rect 152094 0 152150 800
rect 152554 0 152610 800
rect 153014 0 153070 800
rect 153566 0 153622 800
rect 154026 0 154082 800
rect 154486 0 154542 800
rect 154946 0 155002 800
rect 155498 0 155554 800
rect 155958 0 156014 800
rect 156418 0 156474 800
rect 156970 0 157026 800
rect 157430 0 157486 800
rect 157890 0 157946 800
rect 158350 0 158406 800
rect 158902 0 158958 800
rect 159362 0 159418 800
rect 159822 0 159878 800
rect 160374 0 160430 800
rect 160834 0 160890 800
rect 161294 0 161350 800
rect 161754 0 161810 800
rect 162306 0 162362 800
rect 162766 0 162822 800
rect 163226 0 163282 800
rect 163778 0 163834 800
rect 164238 0 164294 800
rect 164698 0 164754 800
rect 165250 0 165306 800
rect 165710 0 165766 800
rect 166170 0 166226 800
rect 166630 0 166686 800
rect 167182 0 167238 800
rect 167642 0 167698 800
rect 168102 0 168158 800
rect 168654 0 168710 800
rect 169114 0 169170 800
rect 169574 0 169630 800
rect 170034 0 170090 800
rect 170586 0 170642 800
rect 171046 0 171102 800
rect 171506 0 171562 800
rect 172058 0 172114 800
rect 172518 0 172574 800
rect 172978 0 173034 800
rect 173438 0 173494 800
rect 173990 0 174046 800
rect 174450 0 174506 800
rect 174910 0 174966 800
rect 175462 0 175518 800
rect 175922 0 175978 800
rect 176382 0 176438 800
rect 176934 0 176990 800
rect 177394 0 177450 800
rect 177854 0 177910 800
rect 178314 0 178370 800
rect 178866 0 178922 800
rect 179326 0 179382 800
rect 179786 0 179842 800
rect 180338 0 180394 800
rect 180798 0 180854 800
rect 181258 0 181314 800
rect 181718 0 181774 800
rect 182270 0 182326 800
rect 182730 0 182786 800
rect 183190 0 183246 800
rect 183742 0 183798 800
rect 184202 0 184258 800
rect 184662 0 184718 800
rect 185122 0 185178 800
rect 185674 0 185730 800
rect 186134 0 186190 800
rect 186594 0 186650 800
rect 187146 0 187202 800
rect 187606 0 187662 800
rect 188066 0 188122 800
rect 188618 0 188674 800
rect 189078 0 189134 800
rect 189538 0 189594 800
rect 189998 0 190054 800
rect 190550 0 190606 800
rect 191010 0 191066 800
rect 191470 0 191526 800
rect 192022 0 192078 800
rect 192482 0 192538 800
rect 192942 0 192998 800
rect 193402 0 193458 800
rect 193954 0 194010 800
rect 194414 0 194470 800
rect 194874 0 194930 800
rect 195426 0 195482 800
rect 195886 0 195942 800
rect 196346 0 196402 800
rect 196898 0 196954 800
rect 197358 0 197414 800
rect 197818 0 197874 800
rect 198278 0 198334 800
rect 198830 0 198886 800
rect 199290 0 199346 800
rect 199750 0 199806 800
rect 200302 0 200358 800
rect 200762 0 200818 800
rect 201222 0 201278 800
rect 201682 0 201738 800
rect 202234 0 202290 800
rect 202694 0 202750 800
rect 203154 0 203210 800
rect 203706 0 203762 800
rect 204166 0 204222 800
rect 204626 0 204682 800
rect 205086 0 205142 800
rect 205638 0 205694 800
rect 206098 0 206154 800
rect 206558 0 206614 800
rect 207110 0 207166 800
rect 207570 0 207626 800
rect 208030 0 208086 800
rect 208582 0 208638 800
rect 209042 0 209098 800
rect 209502 0 209558 800
rect 209962 0 210018 800
rect 210514 0 210570 800
rect 210974 0 211030 800
rect 211434 0 211490 800
rect 211986 0 212042 800
rect 212446 0 212502 800
rect 212906 0 212962 800
rect 213366 0 213422 800
rect 213918 0 213974 800
rect 214378 0 214434 800
rect 214838 0 214894 800
rect 215390 0 215446 800
rect 215850 0 215906 800
rect 216310 0 216366 800
rect 216770 0 216826 800
rect 217322 0 217378 800
rect 217782 0 217838 800
rect 218242 0 218298 800
rect 218794 0 218850 800
rect 219254 0 219310 800
rect 219714 0 219770 800
rect 220266 0 220322 800
rect 220726 0 220782 800
rect 221186 0 221242 800
rect 221646 0 221702 800
rect 222198 0 222254 800
rect 222658 0 222714 800
rect 223118 0 223174 800
rect 223670 0 223726 800
rect 224130 0 224186 800
rect 224590 0 224646 800
rect 225050 0 225106 800
rect 225602 0 225658 800
rect 226062 0 226118 800
rect 226522 0 226578 800
rect 227074 0 227130 800
rect 227534 0 227590 800
rect 227994 0 228050 800
rect 228454 0 228510 800
rect 229006 0 229062 800
rect 229466 0 229522 800
rect 229926 0 229982 800
rect 230478 0 230534 800
rect 230938 0 230994 800
rect 231398 0 231454 800
rect 231950 0 232006 800
rect 232410 0 232466 800
rect 232870 0 232926 800
rect 233330 0 233386 800
rect 233882 0 233938 800
rect 234342 0 234398 800
rect 234802 0 234858 800
rect 235354 0 235410 800
rect 235814 0 235870 800
rect 236274 0 236330 800
rect 236734 0 236790 800
rect 237286 0 237342 800
rect 237746 0 237802 800
rect 238206 0 238262 800
rect 238758 0 238814 800
rect 239218 0 239274 800
rect 239678 0 239734 800
<< obsm2 >>
rect 216 239144 974 239306
rect 1142 239144 2998 239306
rect 3166 239144 5114 239306
rect 5282 239144 7230 239306
rect 7398 239144 9346 239306
rect 9514 239144 11462 239306
rect 11630 239144 13578 239306
rect 13746 239144 15694 239306
rect 15862 239144 17810 239306
rect 17978 239144 19834 239306
rect 20002 239144 21950 239306
rect 22118 239144 24066 239306
rect 24234 239144 26182 239306
rect 26350 239144 28298 239306
rect 28466 239144 30414 239306
rect 30582 239144 32530 239306
rect 32698 239144 34646 239306
rect 34814 239144 36762 239306
rect 36930 239144 38786 239306
rect 38954 239144 40902 239306
rect 41070 239144 43018 239306
rect 43186 239144 45134 239306
rect 45302 239144 47250 239306
rect 47418 239144 49366 239306
rect 49534 239144 51482 239306
rect 51650 239144 53598 239306
rect 53766 239144 55714 239306
rect 55882 239144 57738 239306
rect 57906 239144 59854 239306
rect 60022 239144 61970 239306
rect 62138 239144 64086 239306
rect 64254 239144 66202 239306
rect 66370 239144 68318 239306
rect 68486 239144 70434 239306
rect 70602 239144 72550 239306
rect 72718 239144 74666 239306
rect 74834 239144 76690 239306
rect 76858 239144 78806 239306
rect 78974 239144 80922 239306
rect 81090 239144 83038 239306
rect 83206 239144 85154 239306
rect 85322 239144 87270 239306
rect 87438 239144 89386 239306
rect 89554 239144 91502 239306
rect 91670 239144 93526 239306
rect 93694 239144 95642 239306
rect 95810 239144 97758 239306
rect 97926 239144 99874 239306
rect 100042 239144 101990 239306
rect 102158 239144 104106 239306
rect 104274 239144 106222 239306
rect 106390 239144 108338 239306
rect 108506 239144 110454 239306
rect 110622 239144 112478 239306
rect 112646 239144 114594 239306
rect 114762 239144 116710 239306
rect 116878 239144 118826 239306
rect 118994 239144 120942 239306
rect 121110 239144 123058 239306
rect 123226 239144 125174 239306
rect 125342 239144 127290 239306
rect 127458 239144 129406 239306
rect 129574 239144 131430 239306
rect 131598 239144 133546 239306
rect 133714 239144 135662 239306
rect 135830 239144 137778 239306
rect 137946 239144 139894 239306
rect 140062 239144 142010 239306
rect 142178 239144 144126 239306
rect 144294 239144 146242 239306
rect 146410 239144 148358 239306
rect 148526 239144 150382 239306
rect 150550 239144 152498 239306
rect 152666 239144 154614 239306
rect 154782 239144 156730 239306
rect 156898 239144 158846 239306
rect 159014 239144 160962 239306
rect 161130 239144 163078 239306
rect 163246 239144 165194 239306
rect 165362 239144 167218 239306
rect 167386 239144 169334 239306
rect 169502 239144 171450 239306
rect 171618 239144 173566 239306
rect 173734 239144 175682 239306
rect 175850 239144 177798 239306
rect 177966 239144 179914 239306
rect 180082 239144 182030 239306
rect 182198 239144 184146 239306
rect 184314 239144 186170 239306
rect 186338 239144 188286 239306
rect 188454 239144 190402 239306
rect 190570 239144 192518 239306
rect 192686 239144 194634 239306
rect 194802 239144 196750 239306
rect 196918 239144 198866 239306
rect 199034 239144 200982 239306
rect 201150 239144 203098 239306
rect 203266 239144 205122 239306
rect 205290 239144 207238 239306
rect 207406 239144 209354 239306
rect 209522 239144 211470 239306
rect 211638 239144 213586 239306
rect 213754 239144 215702 239306
rect 215870 239144 217818 239306
rect 217986 239144 219934 239306
rect 220102 239144 222050 239306
rect 222218 239144 224074 239306
rect 224242 239144 226190 239306
rect 226358 239144 228306 239306
rect 228474 239144 230422 239306
rect 230590 239144 232538 239306
rect 232706 239144 234654 239306
rect 234822 239144 236770 239306
rect 236938 239144 238886 239306
rect 239054 239144 239732 239306
rect 216 856 239732 239144
rect 314 2 606 856
rect 774 2 1066 856
rect 1234 2 1526 856
rect 1694 2 2078 856
rect 2246 2 2538 856
rect 2706 2 2998 856
rect 3166 2 3550 856
rect 3718 2 4010 856
rect 4178 2 4470 856
rect 4638 2 4930 856
rect 5098 2 5482 856
rect 5650 2 5942 856
rect 6110 2 6402 856
rect 6570 2 6954 856
rect 7122 2 7414 856
rect 7582 2 7874 856
rect 8042 2 8334 856
rect 8502 2 8886 856
rect 9054 2 9346 856
rect 9514 2 9806 856
rect 9974 2 10358 856
rect 10526 2 10818 856
rect 10986 2 11278 856
rect 11446 2 11830 856
rect 11998 2 12290 856
rect 12458 2 12750 856
rect 12918 2 13210 856
rect 13378 2 13762 856
rect 13930 2 14222 856
rect 14390 2 14682 856
rect 14850 2 15234 856
rect 15402 2 15694 856
rect 15862 2 16154 856
rect 16322 2 16614 856
rect 16782 2 17166 856
rect 17334 2 17626 856
rect 17794 2 18086 856
rect 18254 2 18638 856
rect 18806 2 19098 856
rect 19266 2 19558 856
rect 19726 2 20018 856
rect 20186 2 20570 856
rect 20738 2 21030 856
rect 21198 2 21490 856
rect 21658 2 22042 856
rect 22210 2 22502 856
rect 22670 2 22962 856
rect 23130 2 23514 856
rect 23682 2 23974 856
rect 24142 2 24434 856
rect 24602 2 24894 856
rect 25062 2 25446 856
rect 25614 2 25906 856
rect 26074 2 26366 856
rect 26534 2 26918 856
rect 27086 2 27378 856
rect 27546 2 27838 856
rect 28006 2 28298 856
rect 28466 2 28850 856
rect 29018 2 29310 856
rect 29478 2 29770 856
rect 29938 2 30322 856
rect 30490 2 30782 856
rect 30950 2 31242 856
rect 31410 2 31702 856
rect 31870 2 32254 856
rect 32422 2 32714 856
rect 32882 2 33174 856
rect 33342 2 33726 856
rect 33894 2 34186 856
rect 34354 2 34646 856
rect 34814 2 35198 856
rect 35366 2 35658 856
rect 35826 2 36118 856
rect 36286 2 36578 856
rect 36746 2 37130 856
rect 37298 2 37590 856
rect 37758 2 38050 856
rect 38218 2 38602 856
rect 38770 2 39062 856
rect 39230 2 39522 856
rect 39690 2 39982 856
rect 40150 2 40534 856
rect 40702 2 40994 856
rect 41162 2 41454 856
rect 41622 2 42006 856
rect 42174 2 42466 856
rect 42634 2 42926 856
rect 43094 2 43386 856
rect 43554 2 43938 856
rect 44106 2 44398 856
rect 44566 2 44858 856
rect 45026 2 45410 856
rect 45578 2 45870 856
rect 46038 2 46330 856
rect 46498 2 46882 856
rect 47050 2 47342 856
rect 47510 2 47802 856
rect 47970 2 48262 856
rect 48430 2 48814 856
rect 48982 2 49274 856
rect 49442 2 49734 856
rect 49902 2 50286 856
rect 50454 2 50746 856
rect 50914 2 51206 856
rect 51374 2 51666 856
rect 51834 2 52218 856
rect 52386 2 52678 856
rect 52846 2 53138 856
rect 53306 2 53690 856
rect 53858 2 54150 856
rect 54318 2 54610 856
rect 54778 2 55162 856
rect 55330 2 55622 856
rect 55790 2 56082 856
rect 56250 2 56542 856
rect 56710 2 57094 856
rect 57262 2 57554 856
rect 57722 2 58014 856
rect 58182 2 58566 856
rect 58734 2 59026 856
rect 59194 2 59486 856
rect 59654 2 59946 856
rect 60114 2 60498 856
rect 60666 2 60958 856
rect 61126 2 61418 856
rect 61586 2 61970 856
rect 62138 2 62430 856
rect 62598 2 62890 856
rect 63058 2 63350 856
rect 63518 2 63902 856
rect 64070 2 64362 856
rect 64530 2 64822 856
rect 64990 2 65374 856
rect 65542 2 65834 856
rect 66002 2 66294 856
rect 66462 2 66846 856
rect 67014 2 67306 856
rect 67474 2 67766 856
rect 67934 2 68226 856
rect 68394 2 68778 856
rect 68946 2 69238 856
rect 69406 2 69698 856
rect 69866 2 70250 856
rect 70418 2 70710 856
rect 70878 2 71170 856
rect 71338 2 71630 856
rect 71798 2 72182 856
rect 72350 2 72642 856
rect 72810 2 73102 856
rect 73270 2 73654 856
rect 73822 2 74114 856
rect 74282 2 74574 856
rect 74742 2 75034 856
rect 75202 2 75586 856
rect 75754 2 76046 856
rect 76214 2 76506 856
rect 76674 2 77058 856
rect 77226 2 77518 856
rect 77686 2 77978 856
rect 78146 2 78530 856
rect 78698 2 78990 856
rect 79158 2 79450 856
rect 79618 2 79910 856
rect 80078 2 80462 856
rect 80630 2 80922 856
rect 81090 2 81382 856
rect 81550 2 81934 856
rect 82102 2 82394 856
rect 82562 2 82854 856
rect 83022 2 83314 856
rect 83482 2 83866 856
rect 84034 2 84326 856
rect 84494 2 84786 856
rect 84954 2 85338 856
rect 85506 2 85798 856
rect 85966 2 86258 856
rect 86426 2 86718 856
rect 86886 2 87270 856
rect 87438 2 87730 856
rect 87898 2 88190 856
rect 88358 2 88742 856
rect 88910 2 89202 856
rect 89370 2 89662 856
rect 89830 2 90214 856
rect 90382 2 90674 856
rect 90842 2 91134 856
rect 91302 2 91594 856
rect 91762 2 92146 856
rect 92314 2 92606 856
rect 92774 2 93066 856
rect 93234 2 93618 856
rect 93786 2 94078 856
rect 94246 2 94538 856
rect 94706 2 94998 856
rect 95166 2 95550 856
rect 95718 2 96010 856
rect 96178 2 96470 856
rect 96638 2 97022 856
rect 97190 2 97482 856
rect 97650 2 97942 856
rect 98110 2 98494 856
rect 98662 2 98954 856
rect 99122 2 99414 856
rect 99582 2 99874 856
rect 100042 2 100426 856
rect 100594 2 100886 856
rect 101054 2 101346 856
rect 101514 2 101898 856
rect 102066 2 102358 856
rect 102526 2 102818 856
rect 102986 2 103278 856
rect 103446 2 103830 856
rect 103998 2 104290 856
rect 104458 2 104750 856
rect 104918 2 105302 856
rect 105470 2 105762 856
rect 105930 2 106222 856
rect 106390 2 106682 856
rect 106850 2 107234 856
rect 107402 2 107694 856
rect 107862 2 108154 856
rect 108322 2 108706 856
rect 108874 2 109166 856
rect 109334 2 109626 856
rect 109794 2 110178 856
rect 110346 2 110638 856
rect 110806 2 111098 856
rect 111266 2 111558 856
rect 111726 2 112110 856
rect 112278 2 112570 856
rect 112738 2 113030 856
rect 113198 2 113582 856
rect 113750 2 114042 856
rect 114210 2 114502 856
rect 114670 2 114962 856
rect 115130 2 115514 856
rect 115682 2 115974 856
rect 116142 2 116434 856
rect 116602 2 116986 856
rect 117154 2 117446 856
rect 117614 2 117906 856
rect 118074 2 118366 856
rect 118534 2 118918 856
rect 119086 2 119378 856
rect 119546 2 119838 856
rect 120006 2 120390 856
rect 120558 2 120850 856
rect 121018 2 121310 856
rect 121478 2 121862 856
rect 122030 2 122322 856
rect 122490 2 122782 856
rect 122950 2 123242 856
rect 123410 2 123794 856
rect 123962 2 124254 856
rect 124422 2 124714 856
rect 124882 2 125266 856
rect 125434 2 125726 856
rect 125894 2 126186 856
rect 126354 2 126646 856
rect 126814 2 127198 856
rect 127366 2 127658 856
rect 127826 2 128118 856
rect 128286 2 128670 856
rect 128838 2 129130 856
rect 129298 2 129590 856
rect 129758 2 130050 856
rect 130218 2 130602 856
rect 130770 2 131062 856
rect 131230 2 131522 856
rect 131690 2 132074 856
rect 132242 2 132534 856
rect 132702 2 132994 856
rect 133162 2 133546 856
rect 133714 2 134006 856
rect 134174 2 134466 856
rect 134634 2 134926 856
rect 135094 2 135478 856
rect 135646 2 135938 856
rect 136106 2 136398 856
rect 136566 2 136950 856
rect 137118 2 137410 856
rect 137578 2 137870 856
rect 138038 2 138330 856
rect 138498 2 138882 856
rect 139050 2 139342 856
rect 139510 2 139802 856
rect 139970 2 140354 856
rect 140522 2 140814 856
rect 140982 2 141274 856
rect 141442 2 141734 856
rect 141902 2 142286 856
rect 142454 2 142746 856
rect 142914 2 143206 856
rect 143374 2 143758 856
rect 143926 2 144218 856
rect 144386 2 144678 856
rect 144846 2 145230 856
rect 145398 2 145690 856
rect 145858 2 146150 856
rect 146318 2 146610 856
rect 146778 2 147162 856
rect 147330 2 147622 856
rect 147790 2 148082 856
rect 148250 2 148634 856
rect 148802 2 149094 856
rect 149262 2 149554 856
rect 149722 2 150014 856
rect 150182 2 150566 856
rect 150734 2 151026 856
rect 151194 2 151486 856
rect 151654 2 152038 856
rect 152206 2 152498 856
rect 152666 2 152958 856
rect 153126 2 153510 856
rect 153678 2 153970 856
rect 154138 2 154430 856
rect 154598 2 154890 856
rect 155058 2 155442 856
rect 155610 2 155902 856
rect 156070 2 156362 856
rect 156530 2 156914 856
rect 157082 2 157374 856
rect 157542 2 157834 856
rect 158002 2 158294 856
rect 158462 2 158846 856
rect 159014 2 159306 856
rect 159474 2 159766 856
rect 159934 2 160318 856
rect 160486 2 160778 856
rect 160946 2 161238 856
rect 161406 2 161698 856
rect 161866 2 162250 856
rect 162418 2 162710 856
rect 162878 2 163170 856
rect 163338 2 163722 856
rect 163890 2 164182 856
rect 164350 2 164642 856
rect 164810 2 165194 856
rect 165362 2 165654 856
rect 165822 2 166114 856
rect 166282 2 166574 856
rect 166742 2 167126 856
rect 167294 2 167586 856
rect 167754 2 168046 856
rect 168214 2 168598 856
rect 168766 2 169058 856
rect 169226 2 169518 856
rect 169686 2 169978 856
rect 170146 2 170530 856
rect 170698 2 170990 856
rect 171158 2 171450 856
rect 171618 2 172002 856
rect 172170 2 172462 856
rect 172630 2 172922 856
rect 173090 2 173382 856
rect 173550 2 173934 856
rect 174102 2 174394 856
rect 174562 2 174854 856
rect 175022 2 175406 856
rect 175574 2 175866 856
rect 176034 2 176326 856
rect 176494 2 176878 856
rect 177046 2 177338 856
rect 177506 2 177798 856
rect 177966 2 178258 856
rect 178426 2 178810 856
rect 178978 2 179270 856
rect 179438 2 179730 856
rect 179898 2 180282 856
rect 180450 2 180742 856
rect 180910 2 181202 856
rect 181370 2 181662 856
rect 181830 2 182214 856
rect 182382 2 182674 856
rect 182842 2 183134 856
rect 183302 2 183686 856
rect 183854 2 184146 856
rect 184314 2 184606 856
rect 184774 2 185066 856
rect 185234 2 185618 856
rect 185786 2 186078 856
rect 186246 2 186538 856
rect 186706 2 187090 856
rect 187258 2 187550 856
rect 187718 2 188010 856
rect 188178 2 188562 856
rect 188730 2 189022 856
rect 189190 2 189482 856
rect 189650 2 189942 856
rect 190110 2 190494 856
rect 190662 2 190954 856
rect 191122 2 191414 856
rect 191582 2 191966 856
rect 192134 2 192426 856
rect 192594 2 192886 856
rect 193054 2 193346 856
rect 193514 2 193898 856
rect 194066 2 194358 856
rect 194526 2 194818 856
rect 194986 2 195370 856
rect 195538 2 195830 856
rect 195998 2 196290 856
rect 196458 2 196842 856
rect 197010 2 197302 856
rect 197470 2 197762 856
rect 197930 2 198222 856
rect 198390 2 198774 856
rect 198942 2 199234 856
rect 199402 2 199694 856
rect 199862 2 200246 856
rect 200414 2 200706 856
rect 200874 2 201166 856
rect 201334 2 201626 856
rect 201794 2 202178 856
rect 202346 2 202638 856
rect 202806 2 203098 856
rect 203266 2 203650 856
rect 203818 2 204110 856
rect 204278 2 204570 856
rect 204738 2 205030 856
rect 205198 2 205582 856
rect 205750 2 206042 856
rect 206210 2 206502 856
rect 206670 2 207054 856
rect 207222 2 207514 856
rect 207682 2 207974 856
rect 208142 2 208526 856
rect 208694 2 208986 856
rect 209154 2 209446 856
rect 209614 2 209906 856
rect 210074 2 210458 856
rect 210626 2 210918 856
rect 211086 2 211378 856
rect 211546 2 211930 856
rect 212098 2 212390 856
rect 212558 2 212850 856
rect 213018 2 213310 856
rect 213478 2 213862 856
rect 214030 2 214322 856
rect 214490 2 214782 856
rect 214950 2 215334 856
rect 215502 2 215794 856
rect 215962 2 216254 856
rect 216422 2 216714 856
rect 216882 2 217266 856
rect 217434 2 217726 856
rect 217894 2 218186 856
rect 218354 2 218738 856
rect 218906 2 219198 856
rect 219366 2 219658 856
rect 219826 2 220210 856
rect 220378 2 220670 856
rect 220838 2 221130 856
rect 221298 2 221590 856
rect 221758 2 222142 856
rect 222310 2 222602 856
rect 222770 2 223062 856
rect 223230 2 223614 856
rect 223782 2 224074 856
rect 224242 2 224534 856
rect 224702 2 224994 856
rect 225162 2 225546 856
rect 225714 2 226006 856
rect 226174 2 226466 856
rect 226634 2 227018 856
rect 227186 2 227478 856
rect 227646 2 227938 856
rect 228106 2 228398 856
rect 228566 2 228950 856
rect 229118 2 229410 856
rect 229578 2 229870 856
rect 230038 2 230422 856
rect 230590 2 230882 856
rect 231050 2 231342 856
rect 231510 2 231894 856
rect 232062 2 232354 856
rect 232522 2 232814 856
rect 232982 2 233274 856
rect 233442 2 233826 856
rect 233994 2 234286 856
rect 234454 2 234746 856
rect 234914 2 235298 856
rect 235466 2 235758 856
rect 235926 2 236218 856
rect 236386 2 236678 856
rect 236846 2 237230 856
rect 237398 2 237690 856
rect 237858 2 238150 856
rect 238318 2 238702 856
rect 238870 2 239162 856
rect 239330 2 239622 856
<< obsm3 >>
rect 289 35 234928 237965
<< metal4 >>
rect 4208 2128 4528 237776
rect 19568 2128 19888 237776
rect 34928 2128 35248 237776
rect 50288 2128 50608 237776
rect 65648 2128 65968 237776
rect 81008 2128 81328 237776
rect 96368 2128 96688 237776
rect 111728 2128 112048 237776
rect 127088 2128 127408 237776
rect 142448 2128 142768 237776
rect 157808 2128 158128 237776
rect 173168 2128 173488 237776
rect 188528 2128 188848 237776
rect 203888 2128 204208 237776
rect 219248 2128 219568 237776
rect 234608 2128 234928 237776
<< obsm4 >>
rect 80835 237856 195349 237965
rect 80835 2048 80928 237856
rect 81408 2048 96288 237856
rect 96768 2048 111648 237856
rect 112128 2048 127008 237856
rect 127488 2048 142368 237856
rect 142848 2048 157728 237856
rect 158208 2048 173088 237856
rect 173568 2048 188448 237856
rect 188928 2048 195349 237856
rect 80835 171 195349 2048
<< labels >>
rlabel metal2 s 1030 239200 1086 240000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 64142 239200 64198 240000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 70490 239200 70546 240000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 76746 239200 76802 240000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 83094 239200 83150 240000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 89442 239200 89498 240000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 95698 239200 95754 240000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 102046 239200 102102 240000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 108394 239200 108450 240000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 114650 239200 114706 240000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 120998 239200 121054 240000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 7286 239200 7342 240000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 127346 239200 127402 240000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 133602 239200 133658 240000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 139950 239200 140006 240000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 146298 239200 146354 240000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 152554 239200 152610 240000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 158902 239200 158958 240000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 165250 239200 165306 240000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 171506 239200 171562 240000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 177854 239200 177910 240000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 184202 239200 184258 240000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 13634 239200 13690 240000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 190458 239200 190514 240000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 196806 239200 196862 240000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 203154 239200 203210 240000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 209410 239200 209466 240000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 215758 239200 215814 240000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 222106 239200 222162 240000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 228362 239200 228418 240000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 234710 239200 234766 240000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 19890 239200 19946 240000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 26238 239200 26294 240000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 32586 239200 32642 240000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 38842 239200 38898 240000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 45190 239200 45246 240000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 51538 239200 51594 240000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 57794 239200 57850 240000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3054 239200 3110 240000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 66258 239200 66314 240000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 72606 239200 72662 240000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 78862 239200 78918 240000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 85210 239200 85266 240000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 91558 239200 91614 240000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 97814 239200 97870 240000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 104162 239200 104218 240000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 110510 239200 110566 240000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 116766 239200 116822 240000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 123114 239200 123170 240000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 9402 239200 9458 240000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 129462 239200 129518 240000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 135718 239200 135774 240000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 142066 239200 142122 240000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 148414 239200 148470 240000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 154670 239200 154726 240000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 161018 239200 161074 240000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 167274 239200 167330 240000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 173622 239200 173678 240000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 179970 239200 180026 240000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 186226 239200 186282 240000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 15750 239200 15806 240000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 192574 239200 192630 240000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 198922 239200 198978 240000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 205178 239200 205234 240000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 211526 239200 211582 240000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 217874 239200 217930 240000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 224130 239200 224186 240000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 230478 239200 230534 240000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 236826 239200 236882 240000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 22006 239200 22062 240000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 28354 239200 28410 240000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 34702 239200 34758 240000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 40958 239200 41014 240000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 47306 239200 47362 240000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 53654 239200 53710 240000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 59910 239200 59966 240000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 5170 239200 5226 240000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 68374 239200 68430 240000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 74722 239200 74778 240000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 80978 239200 81034 240000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 87326 239200 87382 240000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 93582 239200 93638 240000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 99930 239200 99986 240000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 106278 239200 106334 240000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 112534 239200 112590 240000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 118882 239200 118938 240000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 125230 239200 125286 240000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 11518 239200 11574 240000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 131486 239200 131542 240000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 137834 239200 137890 240000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 144182 239200 144238 240000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 150438 239200 150494 240000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 156786 239200 156842 240000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 163134 239200 163190 240000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 169390 239200 169446 240000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 175738 239200 175794 240000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 182086 239200 182142 240000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 188342 239200 188398 240000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 17866 239200 17922 240000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 194690 239200 194746 240000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 201038 239200 201094 240000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 207294 239200 207350 240000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 213642 239200 213698 240000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 219990 239200 220046 240000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 226246 239200 226302 240000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 232594 239200 232650 240000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 238942 239200 238998 240000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 24122 239200 24178 240000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 30470 239200 30526 240000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 36818 239200 36874 240000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 43074 239200 43130 240000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 49422 239200 49478 240000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 55770 239200 55826 240000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 62026 239200 62082 240000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 238758 0 238814 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 239218 0 239274 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 239678 0 239734 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 197818 0 197874 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 199290 0 199346 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 200762 0 200818 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 202234 0 202290 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 203706 0 203762 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 205086 0 205142 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 206558 0 206614 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 208030 0 208086 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 209502 0 209558 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 210974 0 211030 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 212446 0 212502 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 213918 0 213974 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 215390 0 215446 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 216770 0 216826 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 218242 0 218298 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 219714 0 219770 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 221186 0 221242 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 222658 0 222714 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 224130 0 224186 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 225602 0 225658 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 227074 0 227130 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 228454 0 228510 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 229926 0 229982 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 231398 0 231454 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 232870 0 232926 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 234342 0 234398 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 235814 0 235870 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 237286 0 237342 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 108762 0 108818 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 123298 0 123354 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 130658 0 130714 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 132130 0 132186 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 134982 0 135038 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 139398 0 139454 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 145286 0 145342 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 146666 0 146722 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 149610 0 149666 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 152554 0 152610 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 154026 0 154082 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 158350 0 158406 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 159822 0 159878 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 161294 0 161350 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 164238 0 164294 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 165710 0 165766 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 167182 0 167238 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 168654 0 168710 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 170034 0 170090 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 171506 0 171562 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 172978 0 173034 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 174450 0 174506 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 175922 0 175978 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 177394 0 177450 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 178866 0 178922 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 180338 0 180394 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 181718 0 181774 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 183190 0 183246 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 184662 0 184718 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 186134 0 186190 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 187606 0 187662 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 189078 0 189134 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 190550 0 190606 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 192022 0 192078 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 193402 0 193458 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 194874 0 194930 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 196346 0 196402 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 198278 0 198334 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 199750 0 199806 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 201222 0 201278 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 202694 0 202750 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 204166 0 204222 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 205638 0 205694 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 207110 0 207166 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 208582 0 208638 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 209962 0 210018 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 211434 0 211490 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 212906 0 212962 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 214378 0 214434 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 215850 0 215906 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 217322 0 217378 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 218794 0 218850 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 220266 0 220322 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 221646 0 221702 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 223118 0 223174 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 224590 0 224646 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 226062 0 226118 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 227534 0 227590 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 229006 0 229062 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 230478 0 230534 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 231950 0 232006 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 233330 0 233386 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 234802 0 234858 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 236274 0 236330 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 237746 0 237802 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 71226 0 71282 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 74170 0 74226 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 77114 0 77170 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 79966 0 80022 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 82910 0 82966 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 85854 0 85910 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 87326 0 87382 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 88798 0 88854 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 90270 0 90326 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 91650 0 91706 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 93122 0 93178 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 94594 0 94650 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 96066 0 96122 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 97538 0 97594 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 99010 0 99066 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 101954 0 102010 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 103334 0 103390 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 104806 0 104862 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 107750 0 107806 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 56598 0 56654 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 110694 0 110750 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 112166 0 112222 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 113638 0 113694 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 115018 0 115074 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 116490 0 116546 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 117962 0 118018 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 119434 0 119490 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 120906 0 120962 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 122378 0 122434 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 123850 0 123906 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 58070 0 58126 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 125322 0 125378 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 126702 0 126758 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 128174 0 128230 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 129646 0 129702 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 131118 0 131174 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 132590 0 132646 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 134062 0 134118 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 135534 0 135590 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 137006 0 137062 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 138386 0 138442 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 139858 0 139914 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 141330 0 141386 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 142802 0 142858 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 144274 0 144330 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 145746 0 145802 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 147218 0 147274 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 148690 0 148746 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 150070 0 150126 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 151542 0 151598 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 153014 0 153070 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 61014 0 61070 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 154486 0 154542 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 155958 0 156014 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 157430 0 157486 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 158902 0 158958 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 161754 0 161810 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 163226 0 163282 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 164698 0 164754 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 166170 0 166226 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 167642 0 167698 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 169114 0 169170 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 170586 0 170642 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 172058 0 172114 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 173438 0 173494 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 174910 0 174966 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 176382 0 176438 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 177854 0 177910 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 179326 0 179382 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 180798 0 180854 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 182270 0 182326 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 183742 0 183798 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 185122 0 185178 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 186594 0 186650 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 188066 0 188122 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 189538 0 189594 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 191010 0 191066 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 192482 0 192538 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 193954 0 194010 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 195426 0 195482 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 196898 0 196954 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 198830 0 198886 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 200302 0 200358 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 201682 0 201738 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 203154 0 203210 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 204626 0 204682 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 206098 0 206154 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 207570 0 207626 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 209042 0 209098 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 210514 0 210570 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 211986 0 212042 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 213366 0 213422 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 214838 0 214894 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 216310 0 216366 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 217782 0 217838 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 219254 0 219310 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 220726 0 220782 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 222198 0 222254 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 223670 0 223726 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 225050 0 225106 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 226522 0 226578 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 227994 0 228050 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 229466 0 229522 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 230938 0 230994 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 232410 0 232466 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 233882 0 233938 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 235354 0 235410 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 236734 0 236790 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 238206 0 238262 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 109682 0 109738 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 111154 0 111210 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 112626 0 112682 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 114098 0 114154 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 119894 0 119950 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 121366 0 121422 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 127254 0 127310 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 134522 0 134578 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 137466 0 137522 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 141790 0 141846 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 143262 0 143318 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 147678 0 147734 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 149150 0 149206 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 150622 0 150678 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 152094 0 152150 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 156418 0 156474 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 157890 0 157946 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 159362 0 159418 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 160834 0 160890 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 162306 0 162362 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 163778 0 163834 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 165250 0 165306 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 166630 0 166686 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 168102 0 168158 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 169574 0 169630 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 171046 0 171102 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 173990 0 174046 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 175462 0 175518 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 176934 0 176990 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 178314 0 178370 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 179786 0 179842 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 181258 0 181314 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 182730 0 182786 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 184202 0 184258 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 185674 0 185730 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 187146 0 187202 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 188618 0 188674 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 191470 0 191526 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 192942 0 192998 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 194414 0 194470 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 195886 0 195942 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 197358 0 197414 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 237776 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 237776 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 237776 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 237776 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 237776 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 237776 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 237776 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 237776 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 237776 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 237776 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 237776 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 237776 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 237776 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 237776 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 237776 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 237776 6 vssd1
port 503 nsew ground input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 662 0 718 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 3054 0 3110 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 36634 0 36690 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 240000 240000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 23790212
string GDS_FILE /root/mar20/tool/caravel_tutorial/caravel_example/openlane/user_proj_example/runs/user_proj_example/results/finishing/user_proj_example.magic.gds
string GDS_START 684714
<< end >>

