magic
tech sky130A
magscale 1 2
timestamp 1647897445
<< metal1 >>
rect 137830 700952 137836 701004
rect 137888 700992 137894 701004
rect 227714 700992 227720 701004
rect 137888 700964 227720 700992
rect 137888 700952 137894 700964
rect 227714 700952 227720 700964
rect 227772 700952 227778 701004
rect 208394 700884 208400 700936
rect 208452 700924 208458 700936
rect 332502 700924 332508 700936
rect 208452 700896 332508 700924
rect 208452 700884 208458 700896
rect 332502 700884 332508 700896
rect 332560 700884 332566 700936
rect 209774 700816 209780 700868
rect 209832 700856 209838 700868
rect 348786 700856 348792 700868
rect 209832 700828 348792 700856
rect 209832 700816 209838 700828
rect 348786 700816 348792 700828
rect 348844 700816 348850 700868
rect 89162 700748 89168 700800
rect 89220 700788 89226 700800
rect 235994 700788 236000 700800
rect 89220 700760 236000 700788
rect 89220 700748 89226 700760
rect 235994 700748 236000 700760
rect 236052 700748 236058 700800
rect 72970 700680 72976 700732
rect 73028 700720 73034 700732
rect 233234 700720 233240 700732
rect 73028 700692 233240 700720
rect 73028 700680 73034 700692
rect 233234 700680 233240 700692
rect 233292 700680 233298 700732
rect 201494 700612 201500 700664
rect 201552 700652 201558 700664
rect 397454 700652 397460 700664
rect 201552 700624 397460 700652
rect 201552 700612 201558 700624
rect 397454 700612 397460 700624
rect 397512 700612 397518 700664
rect 204254 700544 204260 700596
rect 204312 700584 204318 700596
rect 413646 700584 413652 700596
rect 204312 700556 413652 700584
rect 204312 700544 204318 700556
rect 413646 700544 413652 700556
rect 413704 700544 413710 700596
rect 24302 700476 24308 700528
rect 24360 700516 24366 700528
rect 241514 700516 241520 700528
rect 24360 700488 241520 700516
rect 24360 700476 24366 700488
rect 241514 700476 241520 700488
rect 241572 700476 241578 700528
rect 8110 700408 8116 700460
rect 8168 700448 8174 700460
rect 240134 700448 240140 700460
rect 8168 700420 240140 700448
rect 8168 700408 8174 700420
rect 240134 700408 240140 700420
rect 240192 700408 240198 700460
rect 197354 700340 197360 700392
rect 197412 700380 197418 700392
rect 478506 700380 478512 700392
rect 197412 700352 478512 700380
rect 197412 700340 197418 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 191834 700272 191840 700324
rect 191892 700312 191898 700324
rect 543458 700312 543464 700324
rect 191892 700284 543464 700312
rect 191892 700272 191898 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 154114 700204 154120 700256
rect 154172 700244 154178 700256
rect 229094 700244 229100 700256
rect 154172 700216 229100 700244
rect 154172 700204 154178 700216
rect 229094 700204 229100 700216
rect 229152 700204 229158 700256
rect 202782 700136 202788 700188
rect 202840 700176 202846 700188
rect 215938 700176 215944 700188
rect 202840 700148 215944 700176
rect 202840 700136 202846 700148
rect 215938 700136 215944 700148
rect 215996 700136 216002 700188
rect 216674 700136 216680 700188
rect 216732 700176 216738 700188
rect 283834 700176 283840 700188
rect 216732 700148 283840 700176
rect 216732 700136 216738 700148
rect 283834 700136 283840 700148
rect 283892 700136 283898 700188
rect 218974 700068 218980 700120
rect 219032 700108 219038 700120
rect 222194 700108 222200 700120
rect 219032 700080 222200 700108
rect 219032 700068 219038 700080
rect 222194 700068 222200 700080
rect 222252 700068 222258 700120
rect 183554 696940 183560 696992
rect 183612 696980 183618 696992
rect 580166 696980 580172 696992
rect 183612 696952 580172 696980
rect 183612 696940 183618 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 266354 693472 266360 693524
rect 266412 693512 266418 693524
rect 267642 693512 267648 693524
rect 266412 693484 267648 693512
rect 266412 693472 266418 693484
rect 267642 693472 267648 693484
rect 267700 693472 267706 693524
rect 3418 683204 3424 683256
rect 3476 683244 3482 683256
rect 244274 683244 244280 683256
rect 3476 683216 244280 683244
rect 3476 683204 3482 683216
rect 244274 683204 244280 683216
rect 244332 683204 244338 683256
rect 184934 683136 184940 683188
rect 184992 683176 184998 683188
rect 580166 683176 580172 683188
rect 184992 683148 580172 683176
rect 184992 683136 184998 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3418 670760 3424 670812
rect 3476 670800 3482 670812
rect 248414 670800 248420 670812
rect 3476 670772 248420 670800
rect 3476 670760 3482 670772
rect 248414 670760 248420 670772
rect 248472 670760 248478 670812
rect 180794 670692 180800 670744
rect 180852 670732 180858 670744
rect 580166 670732 580172 670744
rect 180852 670704 580172 670732
rect 180852 670692 180858 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 245654 656928 245660 656940
rect 3476 656900 245660 656928
rect 3476 656888 3482 656900
rect 245654 656888 245660 656900
rect 245712 656888 245718 656940
rect 176654 643084 176660 643136
rect 176712 643124 176718 643136
rect 580166 643124 580172 643136
rect 176712 643096 580172 643124
rect 176712 643084 176718 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 249794 632108 249800 632120
rect 3476 632080 249800 632108
rect 3476 632068 3482 632080
rect 249794 632068 249800 632080
rect 249852 632068 249858 632120
rect 178034 630640 178040 630692
rect 178092 630680 178098 630692
rect 580166 630680 580172 630692
rect 178092 630652 580172 630680
rect 178092 630640 178098 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 253934 618304 253940 618316
rect 3200 618276 253940 618304
rect 3200 618264 3206 618276
rect 253934 618264 253940 618276
rect 253992 618264 253998 618316
rect 173894 616836 173900 616888
rect 173952 616876 173958 616888
rect 580166 616876 580172 616888
rect 173952 616848 580172 616876
rect 173952 616836 173958 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 252554 605860 252560 605872
rect 3292 605832 252560 605860
rect 3292 605820 3298 605832
rect 252554 605820 252560 605832
rect 252612 605820 252618 605872
rect 169846 590656 169852 590708
rect 169904 590696 169910 590708
rect 579798 590696 579804 590708
rect 169904 590668 579804 590696
rect 169904 590656 169910 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 256694 579680 256700 579692
rect 3384 579652 256700 579680
rect 3384 579640 3390 579652
rect 256694 579640 256700 579652
rect 256752 579640 256758 579692
rect 172514 576852 172520 576904
rect 172572 576892 172578 576904
rect 580166 576892 580172 576904
rect 172572 576864 580172 576892
rect 172572 576852 172578 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 260834 565876 260840 565888
rect 3476 565848 260840 565876
rect 3476 565836 3482 565848
rect 260834 565836 260840 565848
rect 260892 565836 260898 565888
rect 168374 563048 168380 563100
rect 168432 563088 168438 563100
rect 579798 563088 579804 563100
rect 168432 563060 579804 563088
rect 168432 563048 168438 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 258074 553432 258080 553444
rect 3476 553404 258080 553432
rect 3476 553392 3482 553404
rect 258074 553392 258080 553404
rect 258132 553392 258138 553444
rect 164234 536800 164240 536852
rect 164292 536840 164298 536852
rect 580166 536840 580172 536852
rect 164292 536812 580172 536840
rect 164292 536800 164298 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 262214 527184 262220 527196
rect 3476 527156 262220 527184
rect 3476 527144 3482 527156
rect 262214 527144 262220 527156
rect 262272 527144 262278 527196
rect 165614 524424 165620 524476
rect 165672 524464 165678 524476
rect 580166 524464 580172 524476
rect 165672 524436 580172 524464
rect 165672 524424 165678 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 267734 514808 267740 514820
rect 3476 514780 267740 514808
rect 3476 514768 3482 514780
rect 267734 514768 267740 514780
rect 267792 514768 267798 514820
rect 161474 510620 161480 510672
rect 161532 510660 161538 510672
rect 580166 510660 580172 510672
rect 161532 510632 580172 510660
rect 161532 510620 161538 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 264974 501004 264980 501016
rect 3108 500976 264980 501004
rect 3108 500964 3114 500976
rect 264974 500964 264980 500976
rect 265032 500964 265038 501016
rect 157334 484372 157340 484424
rect 157392 484412 157398 484424
rect 580166 484412 580172 484424
rect 157392 484384 580172 484412
rect 157392 484372 157398 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 269114 474756 269120 474768
rect 3476 474728 269120 474756
rect 3476 474716 3482 474728
rect 269114 474716 269120 474728
rect 269172 474716 269178 474768
rect 160094 470568 160100 470620
rect 160152 470608 160158 470620
rect 579982 470608 579988 470620
rect 160152 470580 579988 470608
rect 160152 470568 160158 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 273254 462380 273260 462392
rect 3292 462352 273260 462380
rect 3292 462340 3298 462352
rect 273254 462340 273260 462352
rect 273312 462340 273318 462392
rect 155954 456764 155960 456816
rect 156012 456804 156018 456816
rect 580166 456804 580172 456816
rect 156012 456776 580172 456804
rect 156012 456764 156018 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 271874 448576 271880 448588
rect 3200 448548 271880 448576
rect 3200 448536 3206 448548
rect 271874 448536 271880 448548
rect 271932 448536 271938 448588
rect 151814 430584 151820 430636
rect 151872 430624 151878 430636
rect 580166 430624 580172 430636
rect 151872 430596 580172 430624
rect 151872 430584 151878 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3418 422288 3424 422340
rect 3476 422328 3482 422340
rect 276014 422328 276020 422340
rect 3476 422300 276020 422328
rect 3476 422288 3482 422300
rect 276014 422288 276020 422300
rect 276072 422288 276078 422340
rect 153194 418140 153200 418192
rect 153252 418180 153258 418192
rect 580166 418180 580172 418192
rect 153252 418152 580172 418180
rect 153252 418140 153258 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 3142 409844 3148 409896
rect 3200 409884 3206 409896
rect 280154 409884 280160 409896
rect 3200 409856 280160 409884
rect 3200 409844 3206 409856
rect 280154 409844 280160 409856
rect 280212 409844 280218 409896
rect 149054 404336 149060 404388
rect 149112 404376 149118 404388
rect 580166 404376 580172 404388
rect 149112 404348 580172 404376
rect 149112 404336 149118 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3418 397468 3424 397520
rect 3476 397508 3482 397520
rect 277394 397508 277400 397520
rect 3476 397480 277400 397508
rect 3476 397468 3482 397480
rect 277394 397468 277400 397480
rect 277452 397468 277458 397520
rect 144914 378156 144920 378208
rect 144972 378196 144978 378208
rect 580166 378196 580172 378208
rect 144972 378168 580172 378196
rect 144972 378156 144978 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 3418 371220 3424 371272
rect 3476 371260 3482 371272
rect 281534 371260 281540 371272
rect 3476 371232 281540 371260
rect 3476 371220 3482 371232
rect 281534 371220 281540 371232
rect 281592 371220 281598 371272
rect 147674 364352 147680 364404
rect 147732 364392 147738 364404
rect 580166 364392 580172 364404
rect 147732 364364 580172 364392
rect 147732 364352 147738 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 284938 357456 284944 357468
rect 3200 357428 284944 357456
rect 3200 357416 3206 357428
rect 284938 357416 284944 357428
rect 284996 357416 285002 357468
rect 143534 351908 143540 351960
rect 143592 351948 143598 351960
rect 580166 351948 580172 351960
rect 143592 351920 580172 351948
rect 143592 351908 143598 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 109402 347760 109408 347812
rect 109460 347800 109466 347812
rect 577682 347800 577688 347812
rect 109460 347772 577688 347800
rect 109460 347760 109466 347772
rect 577682 347760 577688 347772
rect 577740 347760 577746 347812
rect 215110 346332 215116 346384
rect 215168 346372 215174 346384
rect 266354 346372 266360 346384
rect 215168 346344 266360 346372
rect 215168 346332 215174 346344
rect 266354 346332 266360 346344
rect 266412 346332 266418 346384
rect 169754 346264 169760 346316
rect 169812 346304 169818 346316
rect 225598 346304 225604 346316
rect 169812 346276 225604 346304
rect 169812 346264 169818 346276
rect 225598 346264 225604 346276
rect 225656 346264 225662 346316
rect 212994 346196 213000 346248
rect 213052 346236 213058 346248
rect 299474 346236 299480 346248
rect 213052 346208 299480 346236
rect 213052 346196 213058 346208
rect 299474 346196 299480 346208
rect 299532 346196 299538 346248
rect 104894 346128 104900 346180
rect 104952 346168 104958 346180
rect 231946 346168 231952 346180
rect 104952 346140 231952 346168
rect 104952 346128 104958 346140
rect 231946 346128 231952 346140
rect 232004 346128 232010 346180
rect 206646 346060 206652 346112
rect 206704 346100 206710 346112
rect 364334 346100 364340 346112
rect 206704 346072 364340 346100
rect 206704 346060 206710 346072
rect 364334 346060 364340 346072
rect 364392 346060 364398 346112
rect 40034 345992 40040 346044
rect 40092 346032 40098 346044
rect 238294 346032 238300 346044
rect 40092 346004 238300 346032
rect 40092 345992 40098 346004
rect 238294 345992 238300 346004
rect 238352 345992 238358 346044
rect 200390 345924 200396 345976
rect 200448 345964 200454 345976
rect 429194 345964 429200 345976
rect 200448 345936 429200 345964
rect 200448 345924 200454 345936
rect 429194 345924 429200 345936
rect 429252 345924 429258 345976
rect 196158 345856 196164 345908
rect 196216 345896 196222 345908
rect 462314 345896 462320 345908
rect 196216 345868 462320 345896
rect 196216 345856 196222 345868
rect 462314 345856 462320 345868
rect 462372 345856 462378 345908
rect 194042 345788 194048 345840
rect 194100 345828 194106 345840
rect 494054 345828 494060 345840
rect 194100 345800 494060 345828
rect 194100 345788 194106 345800
rect 494054 345788 494060 345800
rect 494112 345788 494118 345840
rect 189810 345720 189816 345772
rect 189868 345760 189874 345772
rect 527174 345760 527180 345772
rect 189868 345732 527180 345760
rect 189868 345720 189874 345732
rect 527174 345720 527180 345732
rect 527232 345720 527238 345772
rect 187694 345652 187700 345704
rect 187752 345692 187758 345704
rect 558914 345692 558920 345704
rect 187752 345664 558920 345692
rect 187752 345652 187758 345664
rect 558914 345652 558920 345664
rect 558972 345652 558978 345704
rect 219342 345584 219348 345636
rect 219400 345624 219406 345636
rect 234614 345624 234620 345636
rect 219400 345596 234620 345624
rect 219400 345584 219406 345596
rect 234614 345584 234620 345596
rect 234672 345584 234678 345636
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 220814 345080 220820 345092
rect 3384 345052 220820 345080
rect 3384 345040 3390 345052
rect 220814 345040 220820 345052
rect 220872 345040 220878 345092
rect 215938 344496 215944 344548
rect 215996 344536 216002 344548
rect 221458 344536 221464 344548
rect 215996 344508 221464 344536
rect 215996 344496 216002 344508
rect 221458 344496 221464 344508
rect 221516 344496 221522 344548
rect 220814 344428 220820 344480
rect 220872 344468 220878 344480
rect 284570 344468 284576 344480
rect 220872 344440 284576 344468
rect 220872 344428 220878 344440
rect 284570 344428 284576 344440
rect 284628 344428 284634 344480
rect 284938 344428 284944 344480
rect 284996 344468 285002 344480
rect 286686 344468 286692 344480
rect 284996 344440 286692 344468
rect 284996 344428 285002 344440
rect 286686 344428 286692 344440
rect 286744 344428 286750 344480
rect 126698 344360 126704 344412
rect 126756 344400 126762 344412
rect 331950 344400 331956 344412
rect 126756 344372 331956 344400
rect 126756 344360 126762 344372
rect 331950 344360 331956 344372
rect 332008 344360 332014 344412
rect 114002 344292 114008 344344
rect 114060 344332 114066 344344
rect 331858 344332 331864 344344
rect 114060 344304 331864 344332
rect 114060 344292 114066 344304
rect 331858 344292 331864 344304
rect 331916 344292 331922 344344
rect 90634 344224 90640 344276
rect 90692 344264 90698 344276
rect 320358 344264 320364 344276
rect 90692 344236 320364 344264
rect 90692 344224 90698 344236
rect 320358 344224 320364 344236
rect 320416 344224 320422 344276
rect 3510 344156 3516 344208
rect 3568 344196 3574 344208
rect 303522 344196 303528 344208
rect 3568 344168 303528 344196
rect 3568 344156 3574 344168
rect 303522 344156 303528 344168
rect 303580 344156 303586 344208
rect 3602 344088 3608 344140
rect 3660 344128 3666 344140
rect 305638 344128 305644 344140
rect 3660 344100 305644 344128
rect 3660 344088 3666 344100
rect 305638 344088 305644 344100
rect 305696 344088 305702 344140
rect 4890 344020 4896 344072
rect 4948 344060 4954 344072
rect 307754 344060 307760 344072
rect 4948 344032 307760 344060
rect 4948 344020 4954 344032
rect 307754 344020 307760 344032
rect 307812 344020 307818 344072
rect 3418 343952 3424 344004
rect 3476 343992 3482 344004
rect 311986 343992 311992 344004
rect 3476 343964 311992 343992
rect 3476 343952 3482 343964
rect 311986 343952 311992 343964
rect 312044 343952 312050 344004
rect 4798 343884 4804 343936
rect 4856 343924 4862 343936
rect 314102 343924 314108 343936
rect 4856 343896 314108 343924
rect 4856 343884 4862 343896
rect 314102 343884 314108 343896
rect 314160 343884 314166 343936
rect 92014 343816 92020 343868
rect 92072 343856 92078 343868
rect 103514 343856 103520 343868
rect 92072 343828 103520 343856
rect 92072 343816 92078 343828
rect 103514 343816 103520 343828
rect 103572 343816 103578 343868
rect 105630 343816 105636 343868
rect 105688 343856 105694 343868
rect 580258 343856 580264 343868
rect 105688 343828 580264 343856
rect 105688 343816 105694 343828
rect 580258 343816 580264 343828
rect 580316 343816 580322 343868
rect 92106 343748 92112 343800
rect 92164 343788 92170 343800
rect 97166 343788 97172 343800
rect 92164 343760 97172 343788
rect 92164 343748 92170 343760
rect 97166 343748 97172 343760
rect 97224 343748 97230 343800
rect 101398 343748 101404 343800
rect 101456 343788 101462 343800
rect 577590 343788 577596 343800
rect 101456 343760 577596 343788
rect 101456 343748 101462 343760
rect 577590 343748 577596 343760
rect 577648 343748 577654 343800
rect 95050 343680 95056 343732
rect 95108 343720 95114 343732
rect 577498 343720 577504 343732
rect 95108 343692 577504 343720
rect 95108 343680 95114 343692
rect 577498 343680 577504 343692
rect 577556 343680 577562 343732
rect 93026 343612 93032 343664
rect 93084 343652 93090 343664
rect 579614 343652 579620 343664
rect 93084 343624 579620 343652
rect 93084 343612 93090 343624
rect 579614 343612 579620 343624
rect 579672 343612 579678 343664
rect 90818 342728 90824 342780
rect 90876 342768 90882 342780
rect 318242 342768 318248 342780
rect 90876 342740 318248 342768
rect 90876 342728 90882 342740
rect 318242 342728 318248 342740
rect 318300 342728 318306 342780
rect 90450 342660 90456 342712
rect 90508 342700 90514 342712
rect 324590 342700 324596 342712
rect 90508 342672 324596 342700
rect 90508 342660 90514 342672
rect 324590 342660 324596 342672
rect 324648 342660 324654 342712
rect 3970 342592 3976 342644
rect 4028 342632 4034 342644
rect 295150 342632 295156 342644
rect 4028 342604 295156 342632
rect 4028 342592 4034 342604
rect 295150 342592 295156 342604
rect 295208 342592 295214 342644
rect 3694 342524 3700 342576
rect 3752 342564 3758 342576
rect 301406 342564 301412 342576
rect 3752 342536 301412 342564
rect 3752 342524 3758 342536
rect 301406 342524 301412 342536
rect 301464 342524 301470 342576
rect 124582 342456 124588 342508
rect 124640 342496 124646 342508
rect 580810 342496 580816 342508
rect 124640 342468 580816 342496
rect 124640 342456 124646 342468
rect 580810 342456 580816 342468
rect 580868 342456 580874 342508
rect 122466 342388 122472 342440
rect 122524 342428 122530 342440
rect 580626 342428 580632 342440
rect 122524 342400 580632 342428
rect 122524 342388 122530 342400
rect 580626 342388 580632 342400
rect 580684 342388 580690 342440
rect 118234 342320 118240 342372
rect 118292 342360 118298 342372
rect 580534 342360 580540 342372
rect 118292 342332 580540 342360
rect 118292 342320 118298 342332
rect 580534 342320 580540 342332
rect 580592 342320 580598 342372
rect 111886 342252 111892 342304
rect 111944 342292 111950 342304
rect 580442 342292 580448 342304
rect 111944 342264 580448 342292
rect 111944 342252 111950 342264
rect 580442 342252 580448 342264
rect 580500 342252 580506 342304
rect 135254 341776 135260 341828
rect 135312 341816 135318 341828
rect 164786 341816 164792 341828
rect 135312 341788 164792 341816
rect 135312 341776 135318 341788
rect 164786 341776 164792 341788
rect 164844 341776 164850 341828
rect 128326 341720 169754 341748
rect 128326 341612 128354 341720
rect 122806 341584 128354 341612
rect 129752 341652 164924 341680
rect 90726 341436 90732 341488
rect 90784 341476 90790 341488
rect 122806 341476 122834 341584
rect 129752 341544 129780 341652
rect 135254 341572 135260 341624
rect 135312 341572 135318 341624
rect 135530 341572 135536 341624
rect 135588 341612 135594 341624
rect 139946 341612 139952 341624
rect 135588 341584 139952 341612
rect 135588 341572 135594 341584
rect 139946 341572 139952 341584
rect 140004 341572 140010 341624
rect 140148 341584 148548 341612
rect 135272 341544 135300 341572
rect 90784 341448 122834 341476
rect 127636 341516 129780 341544
rect 130948 341516 135300 341544
rect 90784 341436 90790 341448
rect 3234 341368 3240 341420
rect 3292 341408 3298 341420
rect 127636 341408 127664 341516
rect 3292 341380 127664 341408
rect 3292 341368 3298 341380
rect 4062 341300 4068 341352
rect 4120 341340 4126 341352
rect 130948 341340 130976 341516
rect 135438 341504 135444 341556
rect 135496 341544 135502 341556
rect 140148 341544 140176 341584
rect 135496 341516 140176 341544
rect 135496 341504 135502 341516
rect 135208 341476 135214 341488
rect 4120 341312 130976 341340
rect 131040 341448 135214 341476
rect 4120 341300 4126 341312
rect 3326 341232 3332 341284
rect 3384 341272 3390 341284
rect 131040 341272 131068 341448
rect 135208 341436 135214 341448
rect 135266 341436 135272 341488
rect 135364 341448 136634 341476
rect 131114 341368 131120 341420
rect 131172 341408 131178 341420
rect 135364 341408 135392 341448
rect 131172 341380 135392 341408
rect 131172 341368 131178 341380
rect 135438 341368 135444 341420
rect 135496 341368 135502 341420
rect 135530 341368 135536 341420
rect 135588 341368 135594 341420
rect 3384 341244 131068 341272
rect 3384 341232 3390 341244
rect 3786 341164 3792 341216
rect 3844 341204 3850 341216
rect 135456 341204 135484 341368
rect 3844 341176 135484 341204
rect 3844 341164 3850 341176
rect 3878 341096 3884 341148
rect 3936 341136 3942 341148
rect 135548 341136 135576 341368
rect 3936 341108 135576 341136
rect 3936 341096 3942 341108
rect 136606 340524 136634 341448
rect 137554 341368 137560 341420
rect 137612 341368 137618 341420
rect 139578 341368 139584 341420
rect 139636 341368 139642 341420
rect 139946 341368 139952 341420
rect 140004 341408 140010 341420
rect 140004 341380 143534 341408
rect 140004 341368 140010 341380
rect 137572 340864 137600 341368
rect 139596 341000 139624 341368
rect 143506 341272 143534 341380
rect 143506 341244 148456 341272
rect 148428 341136 148456 341244
rect 148520 341204 148548 341584
rect 155926 341380 164096 341408
rect 155926 341204 155954 341380
rect 148520 341176 155954 341204
rect 164068 341204 164096 341380
rect 164142 341368 164148 341420
rect 164200 341368 164206 341420
rect 164786 341368 164792 341420
rect 164844 341368 164850 341420
rect 164896 341408 164924 341652
rect 169726 341476 169754 341720
rect 316034 341476 316040 341488
rect 169726 341448 316040 341476
rect 316034 341436 316040 341448
rect 316092 341436 316098 341488
rect 288526 341408 288532 341420
rect 164896 341380 288532 341408
rect 288526 341368 288532 341380
rect 288584 341368 288590 341420
rect 290550 341368 290556 341420
rect 290608 341368 290614 341420
rect 292758 341368 292764 341420
rect 292816 341368 292822 341420
rect 296898 341408 296904 341420
rect 296686 341380 296904 341408
rect 164160 341272 164188 341368
rect 164804 341340 164832 341368
rect 290568 341340 290596 341368
rect 164804 341312 290596 341340
rect 292776 341272 292804 341368
rect 164160 341244 292804 341272
rect 296686 341204 296714 341380
rect 296898 341368 296904 341380
rect 296956 341368 296962 341420
rect 299014 341368 299020 341420
rect 299072 341368 299078 341420
rect 164068 341176 296714 341204
rect 299032 341136 299060 341368
rect 148428 341108 299060 341136
rect 580074 341068 580080 341080
rect 143506 341040 151814 341068
rect 143506 341000 143534 341040
rect 139596 340972 143534 341000
rect 151786 341000 151814 341040
rect 155926 341040 580080 341068
rect 155926 341000 155954 341040
rect 580074 341028 580080 341040
rect 580132 341028 580138 341080
rect 580902 341000 580908 341012
rect 151786 340972 155954 341000
rect 172486 340972 580908 341000
rect 137572 340836 146294 340864
rect 146266 340728 146294 340836
rect 172486 340728 172514 340972
rect 580902 340960 580908 340972
rect 580960 340960 580966 341012
rect 580166 340932 580172 340944
rect 146266 340700 147674 340728
rect 147646 340592 147674 340700
rect 150406 340700 151814 340728
rect 150406 340592 150434 340700
rect 151786 340660 151814 340700
rect 153166 340700 154574 340728
rect 153166 340660 153194 340700
rect 151786 340632 153194 340660
rect 154546 340660 154574 340700
rect 155926 340700 157334 340728
rect 155926 340660 155954 340700
rect 154546 340632 155954 340660
rect 157306 340660 157334 340700
rect 158686 340700 160094 340728
rect 158686 340660 158714 340700
rect 157306 340632 158714 340660
rect 160066 340660 160094 340700
rect 162826 340700 164234 340728
rect 160066 340632 161474 340660
rect 161446 340592 161474 340632
rect 162826 340592 162854 340700
rect 147646 340564 150434 340592
rect 157306 340564 158714 340592
rect 161446 340564 162854 340592
rect 136606 340496 151814 340524
rect 151786 340456 151814 340496
rect 153166 340496 155954 340524
rect 153166 340456 153194 340496
rect 151786 340428 153194 340456
rect 155926 340456 155954 340496
rect 157306 340456 157334 340564
rect 158686 340524 158714 340564
rect 164206 340524 164234 340700
rect 171106 340700 172514 340728
rect 173866 340904 580172 340932
rect 171106 340660 171134 340700
rect 166966 340632 171134 340660
rect 166966 340592 166994 340632
rect 165586 340564 166994 340592
rect 165586 340524 165614 340564
rect 158686 340496 160094 340524
rect 155926 340428 157334 340456
rect 160066 340456 160094 340496
rect 161446 340496 162854 340524
rect 164206 340496 165614 340524
rect 161446 340456 161474 340496
rect 160066 340428 161474 340456
rect 162826 340048 162854 340496
rect 173866 340456 173894 340904
rect 580166 340892 580172 340904
rect 580224 340892 580230 340944
rect 172486 340428 173894 340456
rect 172486 340388 172514 340428
rect 171106 340360 172514 340388
rect 171106 340320 171134 340360
rect 164206 340292 165614 340320
rect 164206 340048 164234 340292
rect 165586 340252 165614 340292
rect 169726 340292 171134 340320
rect 169726 340252 169754 340292
rect 165586 340224 169754 340252
rect 162826 340020 164234 340048
rect 331950 272552 331956 272604
rect 332008 272592 332014 272604
rect 580074 272592 580080 272604
rect 332008 272564 580080 272592
rect 332008 272552 332014 272564
rect 580074 272552 580080 272564
rect 580132 272552 580138 272604
rect 331858 272484 331864 272536
rect 331916 272524 331922 272536
rect 580902 272524 580908 272536
rect 331916 272496 580908 272524
rect 331916 272484 331922 272496
rect 580902 272484 580908 272496
rect 580960 272484 580966 272536
rect 2774 163752 2780 163804
rect 2832 163792 2838 163804
rect 4890 163792 4896 163804
rect 2832 163764 4896 163792
rect 2832 163752 2838 163764
rect 4890 163752 4896 163764
rect 4948 163752 4954 163804
rect 2774 110712 2780 110764
rect 2832 110752 2838 110764
rect 4798 110752 4804 110764
rect 2832 110724 4804 110752
rect 2832 110712 2838 110724
rect 4798 110712 4804 110724
rect 4856 110712 4862 110764
rect 161566 101804 161572 101856
rect 161624 101844 161630 101856
rect 162762 101844 162768 101856
rect 161624 101816 162768 101844
rect 161624 101804 161630 101816
rect 162762 101804 162768 101816
rect 162820 101804 162826 101856
rect 241698 101736 241704 101788
rect 241756 101776 241762 101788
rect 242618 101776 242624 101788
rect 241756 101748 242624 101776
rect 241756 101736 241762 101748
rect 242618 101736 242624 101748
rect 242676 101736 242682 101788
rect 329834 100920 329840 100972
rect 329892 100960 329898 100972
rect 330754 100960 330760 100972
rect 329892 100932 330760 100960
rect 329892 100920 329898 100932
rect 330754 100920 330760 100932
rect 330812 100920 330818 100972
rect 325694 100784 325700 100836
rect 325752 100824 325758 100836
rect 326338 100824 326344 100836
rect 325752 100796 326344 100824
rect 325752 100784 325758 100796
rect 326338 100784 326344 100796
rect 326396 100784 326402 100836
rect 70394 100648 70400 100700
rect 70452 100688 70458 100700
rect 121362 100688 121368 100700
rect 70452 100660 121368 100688
rect 70452 100648 70458 100660
rect 121362 100648 121368 100660
rect 121420 100648 121426 100700
rect 171502 100648 171508 100700
rect 171560 100688 171566 100700
rect 193214 100688 193220 100700
rect 171560 100660 193220 100688
rect 171560 100648 171566 100660
rect 193214 100648 193220 100660
rect 193272 100648 193278 100700
rect 194870 100648 194876 100700
rect 194928 100688 194934 100700
rect 224218 100688 224224 100700
rect 194928 100660 224224 100688
rect 194928 100648 194934 100660
rect 224218 100648 224224 100660
rect 224276 100648 224282 100700
rect 577682 100648 577688 100700
rect 577740 100688 577746 100700
rect 579982 100688 579988 100700
rect 577740 100660 579988 100688
rect 577740 100648 577746 100660
rect 579982 100648 579988 100660
rect 580040 100648 580046 100700
rect 63494 100580 63500 100632
rect 63552 100620 63558 100632
rect 118418 100620 118424 100632
rect 63552 100592 118424 100620
rect 63552 100580 63558 100592
rect 118418 100580 118424 100592
rect 118476 100580 118482 100632
rect 129274 100580 129280 100632
rect 129332 100620 129338 100632
rect 144730 100620 144736 100632
rect 129332 100592 144736 100620
rect 129332 100580 129338 100592
rect 144730 100580 144736 100592
rect 144788 100580 144794 100632
rect 146294 100580 146300 100632
rect 146352 100620 146358 100632
rect 152550 100620 152556 100632
rect 146352 100592 152556 100620
rect 146352 100580 146358 100592
rect 152550 100580 152556 100592
rect 152608 100580 152614 100632
rect 177390 100580 177396 100632
rect 177448 100620 177454 100632
rect 206278 100620 206284 100632
rect 177448 100592 206284 100620
rect 177448 100580 177454 100592
rect 206278 100580 206284 100592
rect 206336 100580 206342 100632
rect 208394 100580 208400 100632
rect 208452 100620 208458 100632
rect 238018 100620 238024 100632
rect 208452 100592 238024 100620
rect 208452 100580 208458 100592
rect 238018 100580 238024 100592
rect 238076 100580 238082 100632
rect 56594 100512 56600 100564
rect 56652 100552 56658 100564
rect 115566 100552 115572 100564
rect 56652 100524 115572 100552
rect 56652 100512 56658 100524
rect 115566 100512 115572 100524
rect 115624 100512 115630 100564
rect 125318 100512 125324 100564
rect 125376 100552 125382 100564
rect 143258 100552 143264 100564
rect 125376 100524 143264 100552
rect 125376 100512 125382 100524
rect 143258 100512 143264 100524
rect 143316 100512 143322 100564
rect 157426 100512 157432 100564
rect 157484 100552 157490 100564
rect 158714 100552 158720 100564
rect 157484 100524 158720 100552
rect 157484 100512 157490 100524
rect 158714 100512 158720 100524
rect 158772 100512 158778 100564
rect 172974 100512 172980 100564
rect 173032 100552 173038 100564
rect 195974 100552 195980 100564
rect 173032 100524 195980 100552
rect 173032 100512 173038 100524
rect 195974 100512 195980 100524
rect 196032 100512 196038 100564
rect 196342 100512 196348 100564
rect 196400 100552 196406 100564
rect 225506 100552 225512 100564
rect 196400 100524 225512 100552
rect 196400 100512 196406 100524
rect 225506 100512 225512 100524
rect 225564 100512 225570 100564
rect 49694 100444 49700 100496
rect 49752 100484 49758 100496
rect 112622 100484 112628 100496
rect 49752 100456 112628 100484
rect 49752 100444 49758 100456
rect 112622 100444 112628 100456
rect 112680 100444 112686 100496
rect 117314 100444 117320 100496
rect 117372 100484 117378 100496
rect 140314 100484 140320 100496
rect 117372 100456 140320 100484
rect 117372 100444 117378 100456
rect 140314 100444 140320 100456
rect 140372 100444 140378 100496
rect 156874 100444 156880 100496
rect 156932 100484 156938 100496
rect 157334 100484 157340 100496
rect 156932 100456 157340 100484
rect 156932 100444 156938 100456
rect 157334 100444 157340 100456
rect 157392 100444 157398 100496
rect 174446 100444 174452 100496
rect 174504 100484 174510 100496
rect 200114 100484 200120 100496
rect 174504 100456 200120 100484
rect 174504 100444 174510 100456
rect 200114 100444 200120 100456
rect 200172 100444 200178 100496
rect 206554 100444 206560 100496
rect 206612 100484 206618 100496
rect 235350 100484 235356 100496
rect 206612 100456 235356 100484
rect 206612 100444 206618 100456
rect 235350 100444 235356 100456
rect 235408 100444 235414 100496
rect 264514 100444 264520 100496
rect 264572 100484 264578 100496
rect 333238 100484 333244 100496
rect 264572 100456 333244 100484
rect 264572 100444 264578 100456
rect 333238 100444 333244 100456
rect 333296 100444 333302 100496
rect 42794 100376 42800 100428
rect 42852 100416 42858 100428
rect 109678 100416 109684 100428
rect 42852 100388 109684 100416
rect 42852 100376 42858 100388
rect 109678 100376 109684 100388
rect 109736 100376 109742 100428
rect 121454 100376 121460 100428
rect 121512 100416 121518 100428
rect 142338 100416 142344 100428
rect 121512 100388 142344 100416
rect 121512 100376 121518 100388
rect 142338 100376 142344 100388
rect 142396 100376 142402 100428
rect 170030 100376 170036 100428
rect 170088 100416 170094 100428
rect 188982 100416 188988 100428
rect 170088 100388 188988 100416
rect 170088 100376 170094 100388
rect 188982 100376 188988 100388
rect 189040 100376 189046 100428
rect 189074 100376 189080 100428
rect 189132 100416 189138 100428
rect 220078 100416 220084 100428
rect 189132 100388 220084 100416
rect 189132 100376 189138 100388
rect 220078 100376 220084 100388
rect 220136 100376 220142 100428
rect 224126 100376 224132 100428
rect 224184 100416 224190 100428
rect 243354 100416 243360 100428
rect 224184 100388 243360 100416
rect 224184 100376 224190 100388
rect 243354 100376 243360 100388
rect 243412 100376 243418 100428
rect 288434 100376 288440 100428
rect 288492 100416 288498 100428
rect 289354 100416 289360 100428
rect 288492 100388 289360 100416
rect 288492 100376 288498 100388
rect 289354 100376 289360 100388
rect 289412 100376 289418 100428
rect 331674 100376 331680 100428
rect 331732 100416 331738 100428
rect 406378 100416 406384 100428
rect 331732 100388 406384 100416
rect 331732 100376 331738 100388
rect 406378 100376 406384 100388
rect 406436 100376 406442 100428
rect 35894 100308 35900 100360
rect 35952 100348 35958 100360
rect 106734 100348 106740 100360
rect 35952 100320 106740 100348
rect 35952 100308 35958 100320
rect 106734 100308 106740 100320
rect 106792 100308 106798 100360
rect 115934 100308 115940 100360
rect 115992 100348 115998 100360
rect 139854 100348 139860 100360
rect 115992 100320 139860 100348
rect 115992 100308 115998 100320
rect 139854 100308 139860 100320
rect 139912 100308 139918 100360
rect 158898 100308 158904 100360
rect 158956 100348 158962 100360
rect 161474 100348 161480 100360
rect 158956 100320 161480 100348
rect 158956 100308 158962 100320
rect 161474 100308 161480 100320
rect 161532 100308 161538 100360
rect 167086 100308 167092 100360
rect 167144 100348 167150 100360
rect 182174 100348 182180 100360
rect 167144 100320 182180 100348
rect 167144 100308 167150 100320
rect 182174 100308 182180 100320
rect 182232 100308 182238 100360
rect 183186 100308 183192 100360
rect 183244 100348 183250 100360
rect 213178 100348 213184 100360
rect 183244 100320 213184 100348
rect 183244 100308 183250 100320
rect 213178 100308 213184 100320
rect 213236 100308 213242 100360
rect 222654 100308 222660 100360
rect 222712 100348 222718 100360
rect 242158 100348 242164 100360
rect 222712 100320 242164 100348
rect 222712 100308 222718 100320
rect 242158 100308 242164 100320
rect 242216 100308 242222 100360
rect 252830 100308 252836 100360
rect 252888 100348 252894 100360
rect 390554 100348 390560 100360
rect 252888 100320 390560 100348
rect 252888 100308 252894 100320
rect 390554 100308 390560 100320
rect 390612 100308 390618 100360
rect 27614 100240 27620 100292
rect 27672 100280 27678 100292
rect 103882 100280 103888 100292
rect 27672 100252 103888 100280
rect 27672 100240 27678 100252
rect 103882 100240 103888 100252
rect 103940 100240 103946 100292
rect 108298 100240 108304 100292
rect 108356 100280 108362 100292
rect 134058 100280 134064 100292
rect 108356 100252 134064 100280
rect 108356 100240 108362 100252
rect 134058 100240 134064 100252
rect 134116 100240 134122 100292
rect 137002 100240 137008 100292
rect 137060 100280 137066 100292
rect 148594 100280 148600 100292
rect 137060 100252 148600 100280
rect 137060 100240 137066 100252
rect 148594 100240 148600 100252
rect 148652 100240 148658 100292
rect 151814 100240 151820 100292
rect 151872 100280 151878 100292
rect 154482 100280 154488 100292
rect 151872 100252 154488 100280
rect 151872 100240 151878 100252
rect 154482 100240 154488 100252
rect 154540 100240 154546 100292
rect 181714 100240 181720 100292
rect 181772 100280 181778 100292
rect 211798 100280 211804 100292
rect 181772 100252 211804 100280
rect 181772 100240 181778 100252
rect 211798 100240 211804 100252
rect 211856 100240 211862 100292
rect 212902 100240 212908 100292
rect 212960 100280 212966 100292
rect 243630 100280 243636 100292
rect 212960 100252 243636 100280
rect 212960 100240 212966 100252
rect 243630 100240 243636 100252
rect 243688 100240 243694 100292
rect 255774 100240 255780 100292
rect 255832 100280 255838 100292
rect 397454 100280 397460 100292
rect 255832 100252 397460 100280
rect 255832 100240 255838 100252
rect 397454 100240 397460 100252
rect 397512 100240 397518 100292
rect 19426 100172 19432 100224
rect 19484 100212 19490 100224
rect 99926 100212 99932 100224
rect 19484 100184 99932 100212
rect 19484 100172 19490 100184
rect 99926 100172 99932 100184
rect 99984 100172 99990 100224
rect 111794 100172 111800 100224
rect 111852 100212 111858 100224
rect 138382 100212 138388 100224
rect 111852 100184 138388 100212
rect 111852 100172 111858 100184
rect 138382 100172 138388 100184
rect 138440 100172 138446 100224
rect 148226 100172 148232 100224
rect 148284 100212 148290 100224
rect 153010 100212 153016 100224
rect 148284 100184 153016 100212
rect 148284 100172 148290 100184
rect 153010 100172 153016 100184
rect 153068 100172 153074 100224
rect 167638 100172 167644 100224
rect 167696 100212 167702 100224
rect 183554 100212 183560 100224
rect 167696 100184 183560 100212
rect 167696 100172 167702 100184
rect 183554 100172 183560 100184
rect 183612 100172 183618 100224
rect 184658 100172 184664 100224
rect 184716 100212 184722 100224
rect 215938 100212 215944 100224
rect 184716 100184 215944 100212
rect 184716 100172 184722 100184
rect 215938 100172 215944 100184
rect 215996 100172 216002 100224
rect 224586 100172 224592 100224
rect 224644 100212 224650 100224
rect 246298 100212 246304 100224
rect 224644 100184 246304 100212
rect 224644 100172 224650 100184
rect 246298 100172 246304 100184
rect 246356 100172 246362 100224
rect 258626 100172 258632 100224
rect 258684 100212 258690 100224
rect 404354 100212 404360 100224
rect 258684 100184 404360 100212
rect 258684 100172 258690 100184
rect 404354 100172 404360 100184
rect 404412 100172 404418 100224
rect 24854 100104 24860 100156
rect 24912 100144 24918 100156
rect 102410 100144 102416 100156
rect 24912 100116 102416 100144
rect 24912 100104 24918 100116
rect 102410 100104 102416 100116
rect 102468 100104 102474 100156
rect 106550 100104 106556 100156
rect 106608 100144 106614 100156
rect 135990 100144 135996 100156
rect 106608 100116 135996 100144
rect 106608 100104 106614 100116
rect 135990 100104 135996 100116
rect 136048 100104 136054 100156
rect 139394 100104 139400 100156
rect 139452 100144 139458 100156
rect 149606 100144 149612 100156
rect 139452 100116 149612 100144
rect 139452 100104 139458 100116
rect 149606 100104 149612 100116
rect 149664 100104 149670 100156
rect 164234 100104 164240 100156
rect 164292 100144 164298 100156
rect 175274 100144 175280 100156
rect 164292 100116 175280 100144
rect 164292 100104 164298 100116
rect 175274 100104 175280 100116
rect 175332 100104 175338 100156
rect 175918 100104 175924 100156
rect 175976 100144 175982 100156
rect 202874 100144 202880 100156
rect 175976 100116 202880 100144
rect 175976 100104 175982 100116
rect 202874 100104 202880 100116
rect 202932 100104 202938 100156
rect 205634 100104 205640 100156
rect 205692 100144 205698 100156
rect 247678 100144 247684 100156
rect 205692 100116 247684 100144
rect 205692 100104 205698 100116
rect 247678 100104 247684 100116
rect 247736 100104 247742 100156
rect 261570 100104 261576 100156
rect 261628 100144 261634 100156
rect 411254 100144 411260 100156
rect 261628 100116 411260 100144
rect 261628 100104 261634 100116
rect 411254 100104 411260 100116
rect 411312 100104 411318 100156
rect 19334 100036 19340 100088
rect 19392 100076 19398 100088
rect 100386 100076 100392 100088
rect 19392 100048 100392 100076
rect 19392 100036 19398 100048
rect 100386 100036 100392 100048
rect 100444 100036 100450 100088
rect 110414 100036 110420 100088
rect 110472 100076 110478 100088
rect 137462 100076 137468 100088
rect 110472 100048 137468 100076
rect 110472 100036 110478 100048
rect 137462 100036 137468 100048
rect 137520 100036 137526 100088
rect 165154 100036 165160 100088
rect 165212 100076 165218 100088
rect 176930 100076 176936 100088
rect 165212 100048 176936 100076
rect 165212 100036 165218 100048
rect 176930 100036 176936 100048
rect 176988 100036 176994 100088
rect 180242 100036 180248 100088
rect 180300 100076 180306 100088
rect 210418 100076 210424 100088
rect 180300 100048 210424 100076
rect 180300 100036 180306 100048
rect 210418 100036 210424 100048
rect 210476 100036 210482 100088
rect 211430 100036 211436 100088
rect 211488 100076 211494 100088
rect 257338 100076 257344 100088
rect 211488 100048 257344 100076
rect 211488 100036 211494 100048
rect 257338 100036 257344 100048
rect 257396 100036 257402 100088
rect 267458 100036 267464 100088
rect 267516 100076 267522 100088
rect 425054 100076 425060 100088
rect 267516 100048 425060 100076
rect 267516 100036 267522 100048
rect 425054 100036 425060 100048
rect 425112 100036 425118 100088
rect 9674 99968 9680 100020
rect 9732 100008 9738 100020
rect 96062 100008 96068 100020
rect 9732 99980 96068 100008
rect 9732 99968 9738 99980
rect 96062 99968 96068 99980
rect 96120 99968 96126 100020
rect 104894 99968 104900 100020
rect 104952 100008 104958 100020
rect 135438 100008 135444 100020
rect 104952 99980 135444 100008
rect 104952 99968 104958 99980
rect 135438 99968 135444 99980
rect 135496 99968 135502 100020
rect 138014 99968 138020 100020
rect 138072 100008 138078 100020
rect 149146 100008 149152 100020
rect 138072 99980 149152 100008
rect 138072 99968 138078 99980
rect 149146 99968 149152 99980
rect 149204 99968 149210 100020
rect 150710 99968 150716 100020
rect 150768 100008 150774 100020
rect 154022 100008 154028 100020
rect 150768 99980 154028 100008
rect 150768 99968 150774 99980
rect 154022 99968 154028 99980
rect 154080 99968 154086 100020
rect 160278 99968 160284 100020
rect 160336 100008 160342 100020
rect 164878 100008 164884 100020
rect 160336 99980 164884 100008
rect 160336 99968 160342 99980
rect 164878 99968 164884 99980
rect 164936 99968 164942 100020
rect 165706 99968 165712 100020
rect 165764 100008 165770 100020
rect 178034 100008 178040 100020
rect 165764 99980 178040 100008
rect 165764 99968 165770 99980
rect 178034 99968 178040 99980
rect 178092 99968 178098 100020
rect 178770 99968 178776 100020
rect 178828 100008 178834 100020
rect 209038 100008 209044 100020
rect 178828 99980 209044 100008
rect 178828 99968 178834 99980
rect 209038 99968 209044 99980
rect 209096 99968 209102 100020
rect 209958 99968 209964 100020
rect 210016 100008 210022 100020
rect 257430 100008 257436 100020
rect 210016 99980 257436 100008
rect 210016 99968 210022 99980
rect 257430 99968 257436 99980
rect 257488 99968 257494 100020
rect 270310 99968 270316 100020
rect 270368 100008 270374 100020
rect 431954 100008 431960 100020
rect 270368 99980 431960 100008
rect 270368 99968 270374 99980
rect 431954 99968 431960 99980
rect 432012 99968 432018 100020
rect 77294 99900 77300 99952
rect 77352 99940 77358 99952
rect 124306 99940 124312 99952
rect 77352 99912 124312 99940
rect 77352 99900 77358 99912
rect 124306 99900 124312 99912
rect 124364 99900 124370 99952
rect 165614 99900 165620 99952
rect 165672 99940 165678 99952
rect 166626 99940 166632 99952
rect 165672 99912 166632 99940
rect 165672 99900 165678 99912
rect 166626 99900 166632 99912
rect 166684 99900 166690 99952
rect 175366 99900 175372 99952
rect 175424 99940 175430 99952
rect 199378 99940 199384 99952
rect 175424 99912 199384 99940
rect 175424 99900 175430 99912
rect 199378 99900 199384 99912
rect 199436 99900 199442 99952
rect 205082 99900 205088 99952
rect 205140 99940 205146 99952
rect 232498 99940 232504 99952
rect 205140 99912 232504 99940
rect 205140 99900 205146 99912
rect 232498 99900 232504 99912
rect 232556 99900 232562 99952
rect 304994 99900 305000 99952
rect 305052 99940 305058 99952
rect 305914 99940 305920 99952
rect 305052 99912 305920 99940
rect 305052 99900 305058 99912
rect 305914 99900 305920 99912
rect 305972 99900 305978 99952
rect 92474 99832 92480 99884
rect 92532 99872 92538 99884
rect 130102 99872 130108 99884
rect 92532 99844 130108 99872
rect 92532 99832 92538 99844
rect 130102 99832 130108 99844
rect 130160 99832 130166 99884
rect 168558 99832 168564 99884
rect 168616 99872 168622 99884
rect 185302 99872 185308 99884
rect 168616 99844 185308 99872
rect 168616 99832 168622 99844
rect 185302 99832 185308 99844
rect 185360 99832 185366 99884
rect 202230 99832 202236 99884
rect 202288 99872 202294 99884
rect 229738 99872 229744 99884
rect 202288 99844 229744 99872
rect 202288 99832 202294 99844
rect 229738 99832 229744 99844
rect 229796 99832 229802 99884
rect 99374 99764 99380 99816
rect 99432 99804 99438 99816
rect 133046 99804 133052 99816
rect 99432 99776 133052 99804
rect 99432 99764 99438 99776
rect 133046 99764 133052 99776
rect 133104 99764 133110 99816
rect 208026 99764 208032 99816
rect 208084 99804 208090 99816
rect 233878 99804 233884 99816
rect 208084 99776 233884 99804
rect 208084 99764 208090 99776
rect 233878 99764 233884 99776
rect 233936 99764 233942 99816
rect 93854 99696 93860 99748
rect 93912 99736 93918 99748
rect 94590 99736 94596 99748
rect 93912 99708 94596 99736
rect 93912 99696 93918 99708
rect 94590 99696 94596 99708
rect 94648 99696 94654 99748
rect 200758 99696 200764 99748
rect 200816 99736 200822 99748
rect 226886 99736 226892 99748
rect 200816 99708 226892 99736
rect 200816 99696 200822 99708
rect 226886 99696 226892 99708
rect 226944 99696 226950 99748
rect 285766 99628 285772 99680
rect 285824 99668 285830 99680
rect 286870 99668 286876 99680
rect 285824 99640 286876 99668
rect 285824 99628 285830 99640
rect 286870 99628 286876 99640
rect 286928 99628 286934 99680
rect 143534 99560 143540 99612
rect 143592 99600 143598 99612
rect 151078 99600 151084 99612
rect 143592 99572 151084 99600
rect 143592 99560 143598 99572
rect 151078 99560 151084 99572
rect 151136 99560 151142 99612
rect 162302 99492 162308 99544
rect 162360 99532 162366 99544
rect 169754 99532 169760 99544
rect 162360 99504 169760 99532
rect 162360 99492 162366 99504
rect 169754 99492 169760 99504
rect 169812 99492 169818 99544
rect 248322 99424 248328 99476
rect 248380 99464 248386 99476
rect 248966 99464 248972 99476
rect 248380 99436 248972 99464
rect 248380 99424 248386 99436
rect 248966 99424 248972 99436
rect 249024 99424 249030 99476
rect 168374 99220 168380 99272
rect 168432 99260 168438 99272
rect 169570 99260 169576 99272
rect 168432 99232 169576 99260
rect 168432 99220 168438 99232
rect 169570 99220 169576 99232
rect 169628 99220 169634 99272
rect 287054 98608 287060 98660
rect 287112 98648 287118 98660
rect 287882 98648 287888 98660
rect 287112 98620 287888 98648
rect 287112 98608 287118 98620
rect 287882 98608 287888 98620
rect 287940 98608 287946 98660
rect 158806 98472 158812 98524
rect 158864 98512 158870 98524
rect 159818 98512 159824 98524
rect 158864 98484 159824 98512
rect 158864 98472 158870 98484
rect 159818 98472 159824 98484
rect 159876 98472 159882 98524
rect 249794 98200 249800 98252
rect 249852 98240 249858 98252
rect 250346 98240 250352 98252
rect 249852 98212 250352 98240
rect 249852 98200 249858 98212
rect 250346 98200 250352 98212
rect 250404 98200 250410 98252
rect 133966 98132 133972 98184
rect 134024 98172 134030 98184
rect 134978 98172 134984 98184
rect 134024 98144 134984 98172
rect 134024 98132 134030 98144
rect 134978 98132 134984 98144
rect 135036 98132 135042 98184
rect 185026 98064 185032 98116
rect 185084 98104 185090 98116
rect 185670 98104 185676 98116
rect 185084 98076 185676 98104
rect 185084 98064 185090 98076
rect 185670 98064 185676 98076
rect 185728 98064 185734 98116
rect 229094 98064 229100 98116
rect 229152 98104 229158 98116
rect 229922 98104 229928 98116
rect 229152 98076 229928 98104
rect 229152 98064 229158 98076
rect 229922 98064 229928 98076
rect 229980 98064 229986 98116
rect 110598 97996 110604 98048
rect 110656 98036 110662 98048
rect 111610 98036 111616 98048
rect 110656 98008 111616 98036
rect 110656 97996 110662 98008
rect 111610 97996 111616 98008
rect 111668 97996 111674 98048
rect 127066 97996 127072 98048
rect 127124 98036 127130 98048
rect 128170 98036 128176 98048
rect 127124 98008 128176 98036
rect 127124 97996 127130 98008
rect 128170 97996 128176 98008
rect 128228 97996 128234 98048
rect 131114 97996 131120 98048
rect 131172 98036 131178 98048
rect 131574 98036 131580 98048
rect 131172 98008 131580 98036
rect 131172 97996 131178 98008
rect 131574 97996 131580 98008
rect 131632 97996 131638 98048
rect 186406 97996 186412 98048
rect 186464 98036 186470 98048
rect 187602 98036 187608 98048
rect 186464 98008 187608 98036
rect 186464 97996 186470 98008
rect 187602 97996 187608 98008
rect 187660 97996 187666 98048
rect 203058 97996 203064 98048
rect 203116 98036 203122 98048
rect 204162 98036 204168 98048
rect 203116 98008 204168 98036
rect 203116 97996 203122 98008
rect 204162 97996 204168 98008
rect 204220 97996 204226 98048
rect 225138 97996 225144 98048
rect 225196 98036 225202 98048
rect 226058 98036 226064 98048
rect 225196 98008 226064 98036
rect 225196 97996 225202 98008
rect 226058 97996 226064 98008
rect 226116 97996 226122 98048
rect 226426 97996 226432 98048
rect 226484 98036 226490 98048
rect 227530 98036 227536 98048
rect 226484 98008 227536 98036
rect 226484 97996 226490 98008
rect 227530 97996 227536 98008
rect 227588 97996 227594 98048
rect 251266 97996 251272 98048
rect 251324 98036 251330 98048
rect 252370 98036 252376 98048
rect 251324 98008 252376 98036
rect 251324 97996 251330 98008
rect 252370 97996 252376 98008
rect 252428 97996 252434 98048
rect 254026 97996 254032 98048
rect 254084 98036 254090 98048
rect 255222 98036 255228 98048
rect 254084 98008 255228 98036
rect 254084 97996 254090 98008
rect 255222 97996 255228 98008
rect 255280 97996 255286 98048
rect 284386 97996 284392 98048
rect 284444 98036 284450 98048
rect 285398 98036 285404 98048
rect 284444 98008 285404 98036
rect 284444 97996 284450 98008
rect 285398 97996 285404 98008
rect 285456 97996 285462 98048
rect 292666 97996 292672 98048
rect 292724 98036 292730 98048
rect 293678 98036 293684 98048
rect 292724 98008 293684 98036
rect 292724 97996 292730 98008
rect 293678 97996 293684 98008
rect 293736 97996 293742 98048
rect 294046 97996 294052 98048
rect 294104 98036 294110 98048
rect 295150 98036 295156 98048
rect 294104 98008 295156 98036
rect 294104 97996 294110 98008
rect 295150 97996 295156 98008
rect 295208 97996 295214 98048
rect 295426 97996 295432 98048
rect 295484 98036 295490 98048
rect 296622 98036 296628 98048
rect 295484 98008 296628 98036
rect 295484 97996 295490 98008
rect 296622 97996 296628 98008
rect 296680 97996 296686 98048
rect 317506 97996 317512 98048
rect 317564 98036 317570 98048
rect 318518 98036 318524 98048
rect 317564 98008 318524 98036
rect 317564 97996 317570 98008
rect 318518 97996 318524 98008
rect 318576 97996 318582 98048
rect 318886 97996 318892 98048
rect 318944 98036 318950 98048
rect 319990 98036 319996 98048
rect 318944 98008 319996 98036
rect 318944 97996 318950 98008
rect 319990 97996 319996 98008
rect 320048 97996 320054 98048
rect 320266 97996 320272 98048
rect 320324 98036 320330 98048
rect 321462 98036 321468 98048
rect 320324 98008 321468 98036
rect 320324 97996 320330 98008
rect 321462 97996 321468 98008
rect 321520 97996 321526 98048
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 90818 97968 90824 97980
rect 3476 97940 90824 97968
rect 3476 97928 3482 97940
rect 90818 97928 90824 97940
rect 90876 97928 90882 97980
rect 91094 97928 91100 97980
rect 91152 97968 91158 97980
rect 92198 97968 92204 97980
rect 91152 97940 92204 97968
rect 91152 97928 91158 97940
rect 92198 97928 92204 97940
rect 92256 97928 92262 97980
rect 92566 97928 92572 97980
rect 92624 97968 92630 97980
rect 93578 97968 93584 97980
rect 92624 97940 93584 97968
rect 92624 97928 92630 97940
rect 93578 97928 93584 97940
rect 93636 97928 93642 97980
rect 100754 97928 100760 97980
rect 100812 97968 100818 97980
rect 101858 97968 101864 97980
rect 100812 97940 101864 97968
rect 100812 97928 100818 97940
rect 101858 97928 101864 97940
rect 101916 97928 101922 97980
rect 102226 97928 102232 97980
rect 102284 97968 102290 97980
rect 103330 97968 103336 97980
rect 102284 97940 103336 97968
rect 102284 97928 102290 97940
rect 103330 97928 103336 97940
rect 103388 97928 103394 97980
rect 103606 97928 103612 97980
rect 103664 97968 103670 97980
rect 104802 97968 104808 97980
rect 103664 97940 104808 97968
rect 103664 97928 103670 97940
rect 104802 97928 104808 97940
rect 104860 97928 104866 97980
rect 107654 97928 107660 97980
rect 107712 97968 107718 97980
rect 108206 97968 108212 97980
rect 107712 97940 108212 97968
rect 107712 97928 107718 97940
rect 108206 97928 108212 97940
rect 108264 97928 108270 97980
rect 110506 97928 110512 97980
rect 110564 97968 110570 97980
rect 111150 97968 111156 97980
rect 110564 97940 111156 97968
rect 110564 97928 110570 97940
rect 111150 97928 111156 97940
rect 111208 97928 111214 97980
rect 113174 97928 113180 97980
rect 113232 97968 113238 97980
rect 114094 97968 114100 97980
rect 113232 97940 114100 97968
rect 113232 97928 113238 97940
rect 114094 97928 114100 97940
rect 114152 97928 114158 97980
rect 118694 97928 118700 97980
rect 118752 97968 118758 97980
rect 119890 97968 119896 97980
rect 118752 97940 119896 97968
rect 118752 97928 118758 97940
rect 119890 97928 119896 97940
rect 119948 97928 119954 97980
rect 120166 97928 120172 97980
rect 120224 97968 120230 97980
rect 120902 97968 120908 97980
rect 120224 97940 120908 97968
rect 120224 97928 120230 97940
rect 120902 97928 120908 97940
rect 120960 97928 120966 97980
rect 126974 97928 126980 97980
rect 127032 97968 127038 97980
rect 127710 97968 127716 97980
rect 127032 97940 127716 97968
rect 127032 97928 127038 97940
rect 127710 97928 127716 97940
rect 127768 97928 127774 97980
rect 131206 97928 131212 97980
rect 131264 97968 131270 97980
rect 132034 97968 132040 97980
rect 131264 97940 132040 97968
rect 131264 97928 131270 97940
rect 132034 97928 132040 97940
rect 132092 97928 132098 97980
rect 140774 97928 140780 97980
rect 140832 97968 140838 97980
rect 141786 97968 141792 97980
rect 140832 97940 141792 97968
rect 140832 97928 140838 97940
rect 141786 97928 141792 97940
rect 141844 97928 141850 97980
rect 143626 97928 143632 97980
rect 143684 97968 143690 97980
rect 144270 97968 144276 97980
rect 143684 97940 144276 97968
rect 143684 97928 143690 97940
rect 144270 97928 144276 97940
rect 144328 97928 144334 97980
rect 144914 97928 144920 97980
rect 144972 97968 144978 97980
rect 145742 97968 145748 97980
rect 144972 97940 145748 97968
rect 144972 97928 144978 97940
rect 145742 97928 145748 97940
rect 145800 97928 145806 97980
rect 146386 97928 146392 97980
rect 146444 97968 146450 97980
rect 147214 97968 147220 97980
rect 146444 97940 147220 97968
rect 146444 97928 146450 97940
rect 147214 97928 147220 97940
rect 147272 97928 147278 97980
rect 160094 97928 160100 97980
rect 160152 97968 160158 97980
rect 161290 97968 161296 97980
rect 160152 97940 161296 97968
rect 160152 97928 160158 97940
rect 161290 97928 161296 97940
rect 161348 97928 161354 97980
rect 169846 97928 169852 97980
rect 169904 97968 169910 97980
rect 171042 97968 171048 97980
rect 169904 97940 171048 97968
rect 169904 97928 169910 97940
rect 171042 97928 171048 97940
rect 171100 97928 171106 97980
rect 178126 97928 178132 97980
rect 178184 97968 178190 97980
rect 179322 97968 179328 97980
rect 178184 97940 179328 97968
rect 178184 97928 178190 97940
rect 179322 97928 179328 97940
rect 179380 97928 179386 97980
rect 185210 97928 185216 97980
rect 185268 97968 185274 97980
rect 186130 97968 186136 97980
rect 185268 97940 186136 97968
rect 185268 97928 185274 97940
rect 186130 97928 186136 97940
rect 186188 97928 186194 97980
rect 186314 97928 186320 97980
rect 186372 97968 186378 97980
rect 187050 97968 187056 97980
rect 186372 97940 187056 97968
rect 186372 97928 186378 97940
rect 187050 97928 187056 97940
rect 187108 97928 187114 97980
rect 189166 97928 189172 97980
rect 189224 97968 189230 97980
rect 189994 97968 190000 97980
rect 189224 97940 190000 97968
rect 189224 97928 189230 97940
rect 189994 97928 190000 97940
rect 190052 97928 190058 97980
rect 190454 97928 190460 97980
rect 190512 97968 190518 97980
rect 191466 97968 191472 97980
rect 190512 97940 191472 97968
rect 190512 97928 190518 97940
rect 191466 97928 191472 97940
rect 191524 97928 191530 97980
rect 191834 97928 191840 97980
rect 191892 97968 191898 97980
rect 192938 97968 192944 97980
rect 191892 97940 192944 97968
rect 191892 97928 191898 97940
rect 192938 97928 192944 97940
rect 192996 97928 193002 97980
rect 194594 97928 194600 97980
rect 194652 97968 194658 97980
rect 195882 97968 195888 97980
rect 194652 97940 195888 97968
rect 194652 97928 194658 97940
rect 195882 97928 195888 97940
rect 195940 97928 195946 97980
rect 202966 97928 202972 97980
rect 203024 97968 203030 97980
rect 203610 97968 203616 97980
rect 203024 97940 203616 97968
rect 203024 97928 203030 97940
rect 203610 97928 203616 97940
rect 203668 97928 203674 97980
rect 208394 97928 208400 97980
rect 208452 97968 208458 97980
rect 209498 97968 209504 97980
rect 208452 97940 209504 97968
rect 208452 97928 208458 97940
rect 209498 97928 209504 97940
rect 209556 97928 209562 97980
rect 209774 97928 209780 97980
rect 209832 97968 209838 97980
rect 210970 97968 210976 97980
rect 209832 97940 210976 97968
rect 209832 97928 209838 97940
rect 210970 97928 210976 97940
rect 211028 97928 211034 97980
rect 211154 97928 211160 97980
rect 211212 97968 211218 97980
rect 212442 97968 212448 97980
rect 211212 97940 212448 97968
rect 211212 97928 211218 97940
rect 212442 97928 212448 97940
rect 212500 97928 212506 97980
rect 224954 97928 224960 97980
rect 225012 97968 225018 97980
rect 225598 97968 225604 97980
rect 225012 97940 225604 97968
rect 225012 97928 225018 97940
rect 225598 97928 225604 97940
rect 225656 97928 225662 97980
rect 226334 97928 226340 97980
rect 226392 97968 226398 97980
rect 226978 97968 226984 97980
rect 226392 97940 226984 97968
rect 226392 97928 226398 97940
rect 226978 97928 226984 97940
rect 227036 97928 227042 97980
rect 227714 97928 227720 97980
rect 227772 97968 227778 97980
rect 228450 97968 228456 97980
rect 227772 97940 228456 97968
rect 227772 97928 227778 97940
rect 228450 97928 228456 97940
rect 228508 97928 228514 97980
rect 230474 97928 230480 97980
rect 230532 97968 230538 97980
rect 231394 97968 231400 97980
rect 230532 97940 231400 97968
rect 230532 97928 230538 97940
rect 231394 97928 231400 97940
rect 231452 97928 231458 97980
rect 233234 97928 233240 97980
rect 233292 97968 233298 97980
rect 234338 97968 234344 97980
rect 233292 97940 234344 97968
rect 233292 97928 233298 97940
rect 234338 97928 234344 97940
rect 234396 97928 234402 97980
rect 234614 97928 234620 97980
rect 234672 97968 234678 97980
rect 235810 97968 235816 97980
rect 234672 97940 235816 97968
rect 234672 97928 234678 97940
rect 235810 97928 235816 97940
rect 235868 97928 235874 97980
rect 241514 97928 241520 97980
rect 241572 97968 241578 97980
rect 242066 97968 242072 97980
rect 241572 97940 242072 97968
rect 241572 97928 241578 97940
rect 242066 97928 242072 97940
rect 242124 97928 242130 97980
rect 242894 97928 242900 97980
rect 242952 97968 242958 97980
rect 243538 97968 243544 97980
rect 242952 97940 243544 97968
rect 242952 97928 242958 97940
rect 243538 97928 243544 97940
rect 243596 97928 243602 97980
rect 244274 97928 244280 97980
rect 244332 97968 244338 97980
rect 245010 97968 245016 97980
rect 244332 97940 245016 97968
rect 244332 97928 244338 97940
rect 245010 97928 245016 97940
rect 245068 97928 245074 97980
rect 248506 97928 248512 97980
rect 248564 97968 248570 97980
rect 249426 97968 249432 97980
rect 248564 97940 249432 97968
rect 248564 97928 248570 97940
rect 249426 97928 249432 97940
rect 249484 97928 249490 97980
rect 251174 97928 251180 97980
rect 251232 97968 251238 97980
rect 251818 97968 251824 97980
rect 251232 97940 251824 97968
rect 251232 97928 251238 97940
rect 251818 97928 251824 97940
rect 251876 97928 251882 97980
rect 253934 97928 253940 97980
rect 253992 97968 253998 97980
rect 254762 97968 254768 97980
rect 253992 97940 254768 97968
rect 253992 97928 253998 97940
rect 254762 97928 254768 97940
rect 254820 97928 254826 97980
rect 258074 97928 258080 97980
rect 258132 97968 258138 97980
rect 259178 97968 259184 97980
rect 258132 97940 259184 97968
rect 258132 97928 258138 97940
rect 259178 97928 259184 97940
rect 259236 97928 259242 97980
rect 259454 97928 259460 97980
rect 259512 97968 259518 97980
rect 260650 97968 260656 97980
rect 259512 97940 260656 97968
rect 259512 97928 259518 97940
rect 260650 97928 260656 97940
rect 260708 97928 260714 97980
rect 260834 97928 260840 97980
rect 260892 97968 260898 97980
rect 262030 97968 262036 97980
rect 260892 97940 262036 97968
rect 260892 97928 260898 97940
rect 262030 97928 262036 97940
rect 262088 97928 262094 97980
rect 262214 97928 262220 97980
rect 262272 97968 262278 97980
rect 263502 97968 263508 97980
rect 262272 97940 263508 97968
rect 262272 97928 262278 97940
rect 263502 97928 263508 97940
rect 263560 97928 263566 97980
rect 266354 97928 266360 97980
rect 266412 97968 266418 97980
rect 266906 97968 266912 97980
rect 266412 97940 266912 97968
rect 266412 97928 266418 97940
rect 266906 97928 266912 97940
rect 266964 97928 266970 97980
rect 267734 97928 267740 97980
rect 267792 97968 267798 97980
rect 268378 97968 268384 97980
rect 267792 97940 268384 97968
rect 267792 97928 267798 97940
rect 268378 97928 268384 97940
rect 268436 97928 268442 97980
rect 269114 97928 269120 97980
rect 269172 97968 269178 97980
rect 269850 97968 269856 97980
rect 269172 97940 269856 97968
rect 269172 97928 269178 97940
rect 269850 97928 269856 97940
rect 269908 97928 269914 97980
rect 270494 97928 270500 97980
rect 270552 97968 270558 97980
rect 271322 97968 271328 97980
rect 270552 97940 271328 97968
rect 270552 97928 270558 97940
rect 271322 97928 271328 97940
rect 271380 97928 271386 97980
rect 271874 97928 271880 97980
rect 271932 97968 271938 97980
rect 272794 97968 272800 97980
rect 271932 97940 272800 97968
rect 271932 97928 271938 97940
rect 272794 97928 272800 97940
rect 272852 97928 272858 97980
rect 282914 97928 282920 97980
rect 282972 97968 282978 97980
rect 283466 97968 283472 97980
rect 282972 97940 283472 97968
rect 282972 97928 282978 97940
rect 283466 97928 283472 97940
rect 283524 97928 283530 97980
rect 284294 97928 284300 97980
rect 284352 97968 284358 97980
rect 284938 97968 284944 97980
rect 284352 97940 284944 97968
rect 284352 97928 284358 97940
rect 284938 97928 284944 97940
rect 284996 97928 285002 97980
rect 285674 97928 285680 97980
rect 285732 97968 285738 97980
rect 286410 97968 286416 97980
rect 285732 97940 286416 97968
rect 285732 97928 285738 97940
rect 286410 97928 286416 97940
rect 286468 97928 286474 97980
rect 287146 97928 287152 97980
rect 287204 97968 287210 97980
rect 288342 97968 288348 97980
rect 287204 97940 288348 97968
rect 287204 97928 287210 97940
rect 288342 97928 288348 97940
rect 288400 97928 288406 97980
rect 291194 97928 291200 97980
rect 291252 97968 291258 97980
rect 291746 97968 291752 97980
rect 291252 97940 291752 97968
rect 291252 97928 291258 97940
rect 291746 97928 291752 97940
rect 291804 97928 291810 97980
rect 292574 97928 292580 97980
rect 292632 97968 292638 97980
rect 293218 97968 293224 97980
rect 292632 97940 293224 97968
rect 292632 97928 292638 97940
rect 293218 97928 293224 97940
rect 293276 97928 293282 97980
rect 293954 97928 293960 97980
rect 294012 97968 294018 97980
rect 294690 97968 294696 97980
rect 294012 97940 294696 97968
rect 294012 97928 294018 97940
rect 294690 97928 294696 97940
rect 294748 97928 294754 97980
rect 295334 97928 295340 97980
rect 295392 97968 295398 97980
rect 296162 97968 296168 97980
rect 295392 97940 296168 97968
rect 295392 97928 295398 97940
rect 296162 97928 296168 97940
rect 296220 97928 296226 97980
rect 299474 97928 299480 97980
rect 299532 97968 299538 97980
rect 300026 97968 300032 97980
rect 299532 97940 300032 97968
rect 299532 97928 299538 97940
rect 300026 97928 300032 97940
rect 300084 97928 300090 97980
rect 300854 97928 300860 97980
rect 300912 97968 300918 97980
rect 301498 97968 301504 97980
rect 300912 97940 301504 97968
rect 300912 97928 300918 97940
rect 301498 97928 301504 97940
rect 301556 97928 301562 97980
rect 302234 97928 302240 97980
rect 302292 97968 302298 97980
rect 302970 97968 302976 97980
rect 302292 97940 302976 97968
rect 302292 97928 302298 97940
rect 302970 97928 302976 97940
rect 303028 97928 303034 97980
rect 303614 97928 303620 97980
rect 303672 97968 303678 97980
rect 304442 97968 304448 97980
rect 303672 97940 304448 97968
rect 303672 97928 303678 97940
rect 304442 97928 304448 97940
rect 304500 97928 304506 97980
rect 307754 97928 307760 97980
rect 307812 97968 307818 97980
rect 308766 97968 308772 97980
rect 307812 97940 308772 97968
rect 307812 97928 307818 97940
rect 308766 97928 308772 97940
rect 308824 97928 308830 97980
rect 309134 97928 309140 97980
rect 309192 97968 309198 97980
rect 310238 97968 310244 97980
rect 309192 97940 310244 97968
rect 309192 97928 309198 97940
rect 310238 97928 310244 97940
rect 310296 97928 310302 97980
rect 310514 97928 310520 97980
rect 310572 97968 310578 97980
rect 311710 97968 311716 97980
rect 310572 97940 311716 97968
rect 310572 97928 310578 97940
rect 311710 97928 311716 97940
rect 311768 97928 311774 97980
rect 311894 97928 311900 97980
rect 311952 97968 311958 97980
rect 313182 97968 313188 97980
rect 311952 97940 313188 97968
rect 311952 97928 311958 97940
rect 313182 97928 313188 97940
rect 313240 97928 313246 97980
rect 317414 97928 317420 97980
rect 317472 97968 317478 97980
rect 318058 97968 318064 97980
rect 317472 97940 318064 97968
rect 317472 97928 317478 97940
rect 318058 97928 318064 97940
rect 318116 97928 318122 97980
rect 318794 97928 318800 97980
rect 318852 97968 318858 97980
rect 319530 97968 319536 97980
rect 318852 97940 319536 97968
rect 318852 97928 318858 97940
rect 319530 97928 319536 97940
rect 319588 97928 319594 97980
rect 320174 97928 320180 97980
rect 320232 97968 320238 97980
rect 321002 97968 321008 97980
rect 320232 97940 321008 97968
rect 320232 97928 320238 97940
rect 321002 97928 321008 97940
rect 321060 97928 321066 97980
rect 321554 97928 321560 97980
rect 321612 97968 321618 97980
rect 322474 97968 322480 97980
rect 321612 97940 322480 97968
rect 321612 97928 321618 97940
rect 322474 97928 322480 97940
rect 322532 97928 322538 97980
rect 324314 97928 324320 97980
rect 324372 97968 324378 97980
rect 324866 97968 324872 97980
rect 324372 97940 324872 97968
rect 324372 97928 324378 97940
rect 324866 97928 324872 97940
rect 324924 97928 324930 97980
rect 327074 97928 327080 97980
rect 327132 97968 327138 97980
rect 327810 97968 327816 97980
rect 327132 97940 327816 97968
rect 327132 97928 327138 97940
rect 327810 97928 327816 97940
rect 327868 97928 327874 97980
rect 328454 97928 328460 97980
rect 328512 97968 328518 97980
rect 329282 97968 329288 97980
rect 328512 97940 329288 97968
rect 328512 97928 328518 97940
rect 329282 97928 329288 97940
rect 329340 97928 329346 97980
rect 92658 97860 92664 97912
rect 92716 97900 92722 97912
rect 93118 97900 93124 97912
rect 92716 97872 93124 97900
rect 92716 97860 92722 97872
rect 93118 97860 93124 97872
rect 93176 97860 93182 97912
rect 97994 97860 98000 97912
rect 98052 97900 98058 97912
rect 98454 97900 98460 97912
rect 98052 97872 98460 97900
rect 98052 97860 98058 97872
rect 98454 97860 98460 97872
rect 98512 97860 98518 97912
rect 116026 97860 116032 97912
rect 116084 97900 116090 97912
rect 116946 97900 116952 97912
rect 116084 97872 116952 97900
rect 116084 97860 116090 97872
rect 116946 97860 116952 97872
rect 117004 97860 117010 97912
rect 136818 97860 136824 97912
rect 136876 97900 136882 97912
rect 137922 97900 137928 97912
rect 136876 97872 137928 97900
rect 136876 97860 136882 97872
rect 137922 97860 137928 97872
rect 137980 97860 137986 97912
rect 140866 97860 140872 97912
rect 140924 97900 140930 97912
rect 141326 97900 141332 97912
rect 140924 97872 141332 97900
rect 140924 97860 140930 97872
rect 141326 97860 141332 97872
rect 141384 97860 141390 97912
rect 176838 97860 176844 97912
rect 176896 97900 176902 97912
rect 177850 97900 177856 97912
rect 176896 97872 177856 97900
rect 176896 97860 176902 97872
rect 177850 97860 177856 97872
rect 177908 97860 177914 97912
rect 197446 97860 197452 97912
rect 197504 97900 197510 97912
rect 198274 97900 198280 97912
rect 197504 97872 198280 97900
rect 197504 97860 197510 97872
rect 198274 97860 198280 97872
rect 198332 97860 198338 97912
rect 198918 97860 198924 97912
rect 198976 97900 198982 97912
rect 199746 97900 199752 97912
rect 198976 97872 199752 97900
rect 198976 97860 198982 97872
rect 199746 97860 199752 97872
rect 199804 97860 199810 97912
rect 215478 97860 215484 97912
rect 215536 97900 215542 97912
rect 216306 97900 216312 97912
rect 215536 97872 216312 97900
rect 215536 97860 215542 97872
rect 216306 97860 216312 97872
rect 216364 97860 216370 97912
rect 216766 97860 216772 97912
rect 216824 97900 216830 97912
rect 217778 97900 217784 97912
rect 216824 97872 217784 97900
rect 216824 97860 216830 97872
rect 217778 97860 217784 97872
rect 217836 97860 217842 97912
rect 218146 97860 218152 97912
rect 218204 97900 218210 97912
rect 219250 97900 219256 97912
rect 218204 97872 219256 97900
rect 218204 97860 218210 97872
rect 219250 97860 219256 97872
rect 219308 97860 219314 97912
rect 220906 97860 220912 97912
rect 220964 97900 220970 97912
rect 222102 97900 222108 97912
rect 220964 97872 222108 97900
rect 220964 97860 220970 97872
rect 222102 97860 222108 97872
rect 222160 97860 222166 97912
rect 229278 97860 229284 97912
rect 229336 97900 229342 97912
rect 230382 97900 230388 97912
rect 229336 97872 230388 97900
rect 229336 97860 229342 97872
rect 230382 97860 230388 97872
rect 230440 97860 230446 97912
rect 231854 97860 231860 97912
rect 231912 97900 231918 97912
rect 232038 97900 232044 97912
rect 231912 97872 232044 97900
rect 231912 97860 231918 97872
rect 232038 97860 232044 97872
rect 232096 97860 232102 97912
rect 237466 97860 237472 97912
rect 237524 97900 237530 97912
rect 238662 97900 238668 97912
rect 237524 97872 238668 97900
rect 237524 97860 237530 97872
rect 238662 97860 238668 97872
rect 238720 97860 238726 97912
rect 249886 97860 249892 97912
rect 249944 97900 249950 97912
rect 250898 97900 250904 97912
rect 249944 97872 250904 97900
rect 249944 97860 249950 97872
rect 250898 97860 250904 97872
rect 250956 97860 250962 97912
rect 256694 97860 256700 97912
rect 256752 97900 256758 97912
rect 257706 97900 257712 97912
rect 256752 97872 257712 97900
rect 256752 97860 256758 97872
rect 257706 97860 257712 97872
rect 257764 97860 257770 97912
rect 289906 97860 289912 97912
rect 289964 97900 289970 97912
rect 290826 97900 290832 97912
rect 289964 97872 290832 97900
rect 289964 97860 289970 97872
rect 290826 97860 290832 97872
rect 290884 97860 290890 97912
rect 291286 97860 291292 97912
rect 291344 97900 291350 97912
rect 292298 97900 292304 97912
rect 291344 97872 292304 97900
rect 291344 97860 291350 97872
rect 292298 97860 292304 97872
rect 292356 97860 292362 97912
rect 298094 97860 298100 97912
rect 298152 97900 298158 97912
rect 298554 97900 298560 97912
rect 298152 97872 298560 97900
rect 298152 97860 298158 97872
rect 298554 97860 298560 97872
rect 298612 97860 298618 97912
rect 306374 97860 306380 97912
rect 306432 97900 306438 97912
rect 307386 97900 307392 97912
rect 306432 97872 307392 97900
rect 306432 97860 306438 97872
rect 307386 97860 307392 97872
rect 307444 97860 307450 97912
rect 323026 97860 323032 97912
rect 323084 97900 323090 97912
rect 323946 97900 323952 97912
rect 323084 97872 323952 97900
rect 323084 97860 323090 97872
rect 323946 97860 323952 97872
rect 324004 97860 324010 97912
rect 324406 97860 324412 97912
rect 324464 97900 324470 97912
rect 325326 97900 325332 97912
rect 324464 97872 325332 97900
rect 324464 97860 324470 97872
rect 325326 97860 325332 97872
rect 325384 97860 325390 97912
rect 106366 97792 106372 97844
rect 106424 97832 106430 97844
rect 107286 97832 107292 97844
rect 106424 97804 107292 97832
rect 106424 97792 106430 97804
rect 107286 97792 107292 97804
rect 107344 97792 107350 97844
rect 107746 97792 107752 97844
rect 107804 97832 107810 97844
rect 108666 97832 108672 97844
rect 107804 97804 108672 97832
rect 107804 97792 107810 97804
rect 108666 97792 108672 97804
rect 108724 97792 108730 97844
rect 180794 97792 180800 97844
rect 180852 97832 180858 97844
rect 181254 97832 181260 97844
rect 180852 97804 181260 97832
rect 180852 97792 180858 97804
rect 181254 97792 181260 97804
rect 181312 97792 181318 97844
rect 182266 97792 182272 97844
rect 182324 97832 182330 97844
rect 182726 97832 182732 97844
rect 182324 97804 182732 97832
rect 182324 97792 182330 97804
rect 182726 97792 182732 97804
rect 182784 97792 182790 97844
rect 183646 97792 183652 97844
rect 183704 97832 183710 97844
rect 184198 97832 184204 97844
rect 183704 97804 184204 97832
rect 183704 97792 183710 97804
rect 184198 97792 184204 97804
rect 184256 97792 184262 97844
rect 197354 97792 197360 97844
rect 197412 97832 197418 97844
rect 197814 97832 197820 97844
rect 197412 97804 197820 97832
rect 197412 97792 197418 97804
rect 197814 97792 197820 97804
rect 197872 97792 197878 97844
rect 200206 97792 200212 97844
rect 200264 97832 200270 97844
rect 201218 97832 201224 97844
rect 200264 97804 201224 97832
rect 200264 97792 200270 97804
rect 201218 97792 201224 97804
rect 201276 97792 201282 97844
rect 240134 97792 240140 97844
rect 240192 97832 240198 97844
rect 240686 97832 240692 97844
rect 240192 97804 240692 97832
rect 240192 97792 240198 97804
rect 240686 97792 240692 97804
rect 240744 97792 240750 97844
rect 243078 97792 243084 97844
rect 243136 97832 243142 97844
rect 244090 97832 244096 97844
rect 243136 97804 244096 97832
rect 243136 97792 243142 97804
rect 244090 97792 244096 97804
rect 244148 97792 244154 97844
rect 281626 97792 281632 97844
rect 281684 97832 281690 97844
rect 282546 97832 282552 97844
rect 281684 97804 282552 97832
rect 281684 97792 281690 97804
rect 282546 97792 282552 97804
rect 282604 97792 282610 97844
rect 283006 97792 283012 97844
rect 283064 97832 283070 97844
rect 284018 97832 284024 97844
rect 283064 97804 284024 97832
rect 283064 97792 283070 97804
rect 284018 97792 284024 97804
rect 284076 97792 284082 97844
rect 289814 97792 289820 97844
rect 289872 97832 289878 97844
rect 290274 97832 290280 97844
rect 289872 97804 290280 97832
rect 289872 97792 289878 97804
rect 290274 97792 290280 97804
rect 290332 97792 290338 97844
rect 322934 97792 322940 97844
rect 322992 97832 322998 97844
rect 323394 97832 323400 97844
rect 322992 97804 323400 97832
rect 322992 97792 322998 97804
rect 323394 97792 323400 97804
rect 323452 97792 323458 97844
rect 128538 97724 128544 97776
rect 128596 97764 128602 97776
rect 129642 97764 129648 97776
rect 128596 97736 129648 97764
rect 128596 97724 128602 97736
rect 129642 97724 129648 97736
rect 129700 97724 129706 97776
rect 219618 97724 219624 97776
rect 219676 97764 219682 97776
rect 220722 97764 220728 97776
rect 219676 97736 220728 97764
rect 219676 97724 219682 97736
rect 220722 97724 220728 97736
rect 220780 97724 220786 97776
rect 231854 97724 231860 97776
rect 231912 97764 231918 97776
rect 232866 97764 232872 97776
rect 231912 97736 232872 97764
rect 231912 97724 231918 97736
rect 232866 97724 232872 97736
rect 232924 97724 232930 97776
rect 245838 97724 245844 97776
rect 245896 97764 245902 97776
rect 246942 97764 246948 97776
rect 245896 97736 246948 97764
rect 245896 97724 245902 97736
rect 246942 97724 246948 97736
rect 247000 97724 247006 97776
rect 281534 97724 281540 97776
rect 281592 97764 281598 97776
rect 281994 97764 282000 97776
rect 281592 97736 282000 97764
rect 281592 97724 281598 97736
rect 281994 97724 282000 97736
rect 282052 97724 282058 97776
rect 106274 96976 106280 97028
rect 106332 97016 106338 97028
rect 106550 97016 106556 97028
rect 106332 96988 106556 97016
rect 106332 96976 106338 96988
rect 106550 96976 106556 96988
rect 106608 96976 106614 97028
rect 147766 94528 147772 94580
rect 147824 94568 147830 94580
rect 148134 94568 148140 94580
rect 147824 94540 148140 94568
rect 147824 94528 147830 94540
rect 148134 94528 148140 94540
rect 148192 94528 148198 94580
rect 150526 94528 150532 94580
rect 150584 94568 150590 94580
rect 151538 94568 151544 94580
rect 150584 94540 151544 94568
rect 150584 94528 150590 94540
rect 151538 94528 151544 94540
rect 151596 94528 151602 94580
rect 154574 94528 154580 94580
rect 154632 94568 154638 94580
rect 155402 94568 155408 94580
rect 154632 94540 155408 94568
rect 154632 94528 154638 94540
rect 155402 94528 155408 94540
rect 155460 94528 155466 94580
rect 155954 94528 155960 94580
rect 156012 94568 156018 94580
rect 156414 94568 156420 94580
rect 156012 94540 156420 94568
rect 156012 94528 156018 94540
rect 156414 94528 156420 94540
rect 156472 94528 156478 94580
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 90726 85524 90732 85536
rect 3200 85496 90732 85524
rect 3200 85484 3206 85496
rect 90726 85484 90732 85496
rect 90784 85484 90790 85536
rect 577590 73108 577596 73160
rect 577648 73148 577654 73160
rect 579706 73148 579712 73160
rect 577648 73120 579712 73148
rect 577648 73108 577654 73120
rect 579706 73108 579712 73120
rect 579764 73108 579770 73160
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 90634 71720 90640 71732
rect 3476 71692 90640 71720
rect 3476 71680 3482 71692
rect 90634 71680 90640 71692
rect 90692 71680 90698 71732
rect 92014 60664 92020 60716
rect 92072 60704 92078 60716
rect 580166 60704 580172 60716
rect 92072 60676 580172 60704
rect 92072 60664 92078 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 90450 59344 90456 59356
rect 3108 59316 90456 59344
rect 3108 59304 3114 59316
rect 90450 59304 90456 59316
rect 90508 59304 90514 59356
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 90542 45540 90548 45552
rect 3476 45512 90548 45540
rect 3476 45500 3482 45512
rect 90542 45500 90548 45512
rect 90600 45500 90606 45552
rect 3142 33056 3148 33108
rect 3200 33096 3206 33108
rect 90358 33096 90364 33108
rect 3200 33068 90364 33096
rect 3200 33056 3206 33068
rect 90358 33056 90364 33068
rect 90416 33056 90422 33108
rect 577498 33056 577504 33108
rect 577556 33096 577562 33108
rect 579614 33096 579620 33108
rect 577556 33068 579620 33096
rect 577556 33056 577562 33068
rect 579614 33056 579620 33068
rect 579672 33056 579678 33108
rect 254118 23128 254124 23180
rect 254176 23168 254182 23180
rect 393314 23168 393320 23180
rect 254176 23140 393320 23168
rect 254176 23128 254182 23140
rect 393314 23128 393320 23140
rect 393372 23128 393378 23180
rect 256878 23060 256884 23112
rect 256936 23100 256942 23112
rect 400214 23100 400220 23112
rect 256936 23072 400220 23100
rect 256936 23060 256942 23072
rect 400214 23060 400220 23072
rect 400272 23060 400278 23112
rect 259638 22992 259644 23044
rect 259696 23032 259702 23044
rect 407114 23032 407120 23044
rect 259696 23004 407120 23032
rect 259696 22992 259702 23004
rect 407114 22992 407120 23004
rect 407172 22992 407178 23044
rect 262398 22924 262404 22976
rect 262456 22964 262462 22976
rect 415394 22964 415400 22976
rect 262456 22936 415400 22964
rect 262456 22924 262462 22936
rect 415394 22924 415400 22936
rect 415452 22924 415458 22976
rect 265158 22856 265164 22908
rect 265216 22896 265222 22908
rect 422294 22896 422300 22908
rect 265216 22868 422300 22896
rect 265216 22856 265222 22868
rect 422294 22856 422300 22868
rect 422352 22856 422358 22908
rect 267918 22788 267924 22840
rect 267976 22828 267982 22840
rect 429194 22828 429200 22840
rect 267976 22800 429200 22828
rect 267976 22788 267982 22800
rect 429194 22788 429200 22800
rect 429252 22788 429258 22840
rect 270678 22720 270684 22772
rect 270736 22760 270742 22772
rect 436094 22760 436100 22772
rect 270736 22732 436100 22760
rect 270736 22720 270742 22732
rect 436094 22720 436100 22732
rect 436152 22720 436158 22772
rect 240318 22040 240324 22092
rect 240376 22080 240382 22092
rect 361574 22080 361580 22092
rect 240376 22052 361580 22080
rect 240376 22040 240382 22052
rect 361574 22040 361580 22052
rect 361632 22040 361638 22092
rect 241698 21972 241704 22024
rect 241756 22012 241762 22024
rect 365714 22012 365720 22024
rect 241756 21984 365720 22012
rect 241756 21972 241762 21984
rect 365714 21972 365720 21984
rect 365772 21972 365778 22024
rect 243078 21904 243084 21956
rect 243136 21944 243142 21956
rect 368474 21944 368480 21956
rect 243136 21916 368480 21944
rect 243136 21904 243142 21916
rect 368474 21904 368480 21916
rect 368532 21904 368538 21956
rect 244458 21836 244464 21888
rect 244516 21876 244522 21888
rect 372614 21876 372620 21888
rect 244516 21848 372620 21876
rect 244516 21836 244522 21848
rect 372614 21836 372620 21848
rect 372672 21836 372678 21888
rect 245838 21768 245844 21820
rect 245896 21808 245902 21820
rect 375374 21808 375380 21820
rect 245896 21780 375380 21808
rect 245896 21768 245902 21780
rect 375374 21768 375380 21780
rect 375432 21768 375438 21820
rect 248598 21700 248604 21752
rect 248656 21740 248662 21752
rect 379514 21740 379520 21752
rect 248656 21712 379520 21740
rect 248656 21700 248662 21712
rect 379514 21700 379520 21712
rect 379572 21700 379578 21752
rect 249978 21632 249984 21684
rect 250036 21672 250042 21684
rect 382274 21672 382280 21684
rect 250036 21644 382280 21672
rect 250036 21632 250042 21644
rect 382274 21632 382280 21644
rect 382332 21632 382338 21684
rect 251358 21564 251364 21616
rect 251416 21604 251422 21616
rect 386414 21604 386420 21616
rect 251416 21576 386420 21604
rect 251416 21564 251422 21576
rect 386414 21564 386420 21576
rect 386472 21564 386478 21616
rect 309318 21496 309324 21548
rect 309376 21536 309382 21548
rect 528554 21536 528560 21548
rect 309376 21508 528560 21536
rect 309376 21496 309382 21508
rect 528554 21496 528560 21508
rect 528612 21496 528618 21548
rect 310698 21428 310704 21480
rect 310756 21468 310762 21480
rect 531314 21468 531320 21480
rect 310756 21440 531320 21468
rect 310756 21428 310762 21440
rect 531314 21428 531320 21440
rect 531372 21428 531378 21480
rect 312078 21360 312084 21412
rect 312136 21400 312142 21412
rect 535454 21400 535460 21412
rect 312136 21372 535460 21400
rect 312136 21360 312142 21372
rect 535454 21360 535460 21372
rect 535512 21360 535518 21412
rect 238846 21292 238852 21344
rect 238904 21332 238910 21344
rect 357434 21332 357440 21344
rect 238904 21304 357440 21332
rect 238904 21292 238910 21304
rect 357434 21292 357440 21304
rect 357492 21292 357498 21344
rect 237558 21224 237564 21276
rect 237616 21264 237622 21276
rect 354674 21264 354680 21276
rect 237616 21236 354680 21264
rect 237616 21224 237622 21236
rect 354674 21224 354680 21236
rect 354732 21224 354738 21276
rect 236178 21156 236184 21208
rect 236236 21196 236242 21208
rect 350534 21196 350540 21208
rect 236236 21168 350540 21196
rect 236236 21156 236242 21168
rect 350534 21156 350540 21168
rect 350592 21156 350598 21208
rect 92106 20612 92112 20664
rect 92164 20652 92170 20664
rect 579982 20652 579988 20664
rect 92164 20624 579988 20652
rect 92164 20612 92170 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 252646 20544 252652 20596
rect 252704 20584 252710 20596
rect 391934 20584 391940 20596
rect 252704 20556 391940 20584
rect 252704 20544 252710 20556
rect 391934 20544 391940 20556
rect 391992 20544 391998 20596
rect 254026 20476 254032 20528
rect 254084 20516 254090 20528
rect 396074 20516 396080 20528
rect 254084 20488 396080 20516
rect 254084 20476 254090 20488
rect 396074 20476 396080 20488
rect 396132 20476 396138 20528
rect 256786 20408 256792 20460
rect 256844 20448 256850 20460
rect 398834 20448 398840 20460
rect 256844 20420 398840 20448
rect 256844 20408 256850 20420
rect 398834 20408 398840 20420
rect 398892 20408 398898 20460
rect 258166 20340 258172 20392
rect 258224 20380 258230 20392
rect 402974 20380 402980 20392
rect 258224 20352 402980 20380
rect 258224 20340 258230 20352
rect 402974 20340 402980 20352
rect 403032 20340 403038 20392
rect 278958 20272 278964 20324
rect 279016 20312 279022 20324
rect 456886 20312 456892 20324
rect 279016 20284 456892 20312
rect 279016 20272 279022 20284
rect 456886 20272 456892 20284
rect 456944 20272 456950 20324
rect 281718 20204 281724 20256
rect 281776 20244 281782 20256
rect 459554 20244 459560 20256
rect 281776 20216 459560 20244
rect 281776 20204 281782 20216
rect 459554 20204 459560 20216
rect 459612 20204 459618 20256
rect 283098 20136 283104 20188
rect 283156 20176 283162 20188
rect 463694 20176 463700 20188
rect 283156 20148 463700 20176
rect 283156 20136 283162 20148
rect 463694 20136 463700 20148
rect 463752 20136 463758 20188
rect 284478 20068 284484 20120
rect 284536 20108 284542 20120
rect 466454 20108 466460 20120
rect 284536 20080 466460 20108
rect 284536 20068 284542 20080
rect 466454 20068 466460 20080
rect 466512 20068 466518 20120
rect 285858 20000 285864 20052
rect 285916 20040 285922 20052
rect 470594 20040 470600 20052
rect 285916 20012 470600 20040
rect 285916 20000 285922 20012
rect 470594 20000 470600 20012
rect 470652 20000 470658 20052
rect 307938 19932 307944 19984
rect 307996 19972 308002 19984
rect 524414 19972 524420 19984
rect 307996 19944 524420 19972
rect 307996 19932 308002 19944
rect 524414 19932 524420 19944
rect 524472 19932 524478 19984
rect 251266 19864 251272 19916
rect 251324 19904 251330 19916
rect 389174 19904 389180 19916
rect 251324 19876 389180 19904
rect 251324 19864 251330 19876
rect 389174 19864 389180 19876
rect 389232 19864 389238 19916
rect 234798 19796 234804 19848
rect 234856 19836 234862 19848
rect 347774 19836 347780 19848
rect 234856 19808 347780 19836
rect 234856 19796 234862 19808
rect 347774 19796 347780 19808
rect 347832 19796 347838 19848
rect 232038 19728 232044 19780
rect 232096 19768 232102 19780
rect 339494 19768 339500 19780
rect 232096 19740 339500 19768
rect 232096 19728 232102 19740
rect 339494 19728 339500 19740
rect 339552 19728 339558 19780
rect 267826 19252 267832 19304
rect 267884 19292 267890 19304
rect 426434 19292 426440 19304
rect 267884 19264 426440 19292
rect 267884 19252 267890 19264
rect 426434 19252 426440 19264
rect 426492 19252 426498 19304
rect 269206 19184 269212 19236
rect 269264 19224 269270 19236
rect 430574 19224 430580 19236
rect 269264 19196 430580 19224
rect 269264 19184 269270 19196
rect 430574 19184 430580 19196
rect 430632 19184 430638 19236
rect 270586 19116 270592 19168
rect 270644 19156 270650 19168
rect 433334 19156 433340 19168
rect 270644 19128 433340 19156
rect 270644 19116 270650 19128
rect 433334 19116 433340 19128
rect 433392 19116 433398 19168
rect 271966 19048 271972 19100
rect 272024 19088 272030 19100
rect 437474 19088 437480 19100
rect 272024 19060 437480 19088
rect 272024 19048 272030 19060
rect 437474 19048 437480 19060
rect 437532 19048 437538 19100
rect 298278 18980 298284 19032
rect 298336 19020 298342 19032
rect 502334 19020 502340 19032
rect 298336 18992 502340 19020
rect 298336 18980 298342 18992
rect 502334 18980 502340 18992
rect 502392 18980 502398 19032
rect 299658 18912 299664 18964
rect 299716 18952 299722 18964
rect 506474 18952 506480 18964
rect 299716 18924 506480 18952
rect 299716 18912 299722 18924
rect 506474 18912 506480 18924
rect 506532 18912 506538 18964
rect 301038 18844 301044 18896
rect 301096 18884 301102 18896
rect 509234 18884 509240 18896
rect 301096 18856 509240 18884
rect 301096 18844 301102 18856
rect 509234 18844 509240 18856
rect 509292 18844 509298 18896
rect 302418 18776 302424 18828
rect 302476 18816 302482 18828
rect 513374 18816 513380 18828
rect 302476 18788 513380 18816
rect 302476 18776 302482 18788
rect 513374 18776 513380 18788
rect 513432 18776 513438 18828
rect 303798 18708 303804 18760
rect 303856 18748 303862 18760
rect 516134 18748 516140 18760
rect 303856 18720 516140 18748
rect 303856 18708 303862 18720
rect 516134 18708 516140 18720
rect 516192 18708 516198 18760
rect 325878 18640 325884 18692
rect 325936 18680 325942 18692
rect 569954 18680 569960 18692
rect 325936 18652 569960 18680
rect 325936 18640 325942 18652
rect 569954 18640 569960 18652
rect 570012 18640 570018 18692
rect 327258 18572 327264 18624
rect 327316 18612 327322 18624
rect 572714 18612 572720 18624
rect 327316 18584 572720 18612
rect 327316 18572 327322 18584
rect 572714 18572 572720 18584
rect 572772 18572 572778 18624
rect 266446 18504 266452 18556
rect 266504 18544 266510 18556
rect 423674 18544 423680 18556
rect 266504 18516 423680 18544
rect 266504 18504 266510 18516
rect 423674 18504 423680 18516
rect 423732 18504 423738 18556
rect 229278 18436 229284 18488
rect 229336 18476 229342 18488
rect 335354 18476 335360 18488
rect 229336 18448 335360 18476
rect 229336 18436 229342 18448
rect 335354 18436 335360 18448
rect 335412 18436 335418 18488
rect 227898 18368 227904 18420
rect 227956 18408 227962 18420
rect 332594 18408 332600 18420
rect 227956 18380 332600 18408
rect 227956 18368 227962 18380
rect 332594 18368 332600 18380
rect 332652 18368 332658 18420
rect 242986 17892 242992 17944
rect 243044 17932 243050 17944
rect 365806 17932 365812 17944
rect 243044 17904 365812 17932
rect 243044 17892 243050 17904
rect 365806 17892 365812 17904
rect 365864 17892 365870 17944
rect 244366 17824 244372 17876
rect 244424 17864 244430 17876
rect 369854 17864 369860 17876
rect 244424 17836 369860 17864
rect 244424 17824 244430 17836
rect 369854 17824 369860 17836
rect 369912 17824 369918 17876
rect 289998 17756 290004 17808
rect 290056 17796 290062 17808
rect 480254 17796 480260 17808
rect 290056 17768 480260 17796
rect 290056 17756 290062 17768
rect 480254 17756 480260 17768
rect 480312 17756 480318 17808
rect 291378 17688 291384 17740
rect 291436 17728 291442 17740
rect 483014 17728 483020 17740
rect 291436 17700 483020 17728
rect 291436 17688 291442 17700
rect 483014 17688 483020 17700
rect 483072 17688 483078 17740
rect 292758 17620 292764 17672
rect 292816 17660 292822 17672
rect 487154 17660 487160 17672
rect 292816 17632 487160 17660
rect 292816 17620 292822 17632
rect 487154 17620 487160 17632
rect 487212 17620 487218 17672
rect 294138 17552 294144 17604
rect 294196 17592 294202 17604
rect 489914 17592 489920 17604
rect 294196 17564 489920 17592
rect 294196 17552 294202 17564
rect 489914 17552 489920 17564
rect 489972 17552 489978 17604
rect 295518 17484 295524 17536
rect 295576 17524 295582 17536
rect 494054 17524 494060 17536
rect 295576 17496 494060 17524
rect 295576 17484 295582 17496
rect 494054 17484 494060 17496
rect 494112 17484 494118 17536
rect 317598 17416 317604 17468
rect 317656 17456 317662 17468
rect 547874 17456 547880 17468
rect 317656 17428 547880 17456
rect 317656 17416 317662 17428
rect 547874 17416 547880 17428
rect 547932 17416 547938 17468
rect 318978 17348 318984 17400
rect 319036 17388 319042 17400
rect 550634 17388 550640 17400
rect 319036 17360 550640 17388
rect 319036 17348 319042 17360
rect 550634 17348 550640 17360
rect 550692 17348 550698 17400
rect 320358 17280 320364 17332
rect 320416 17320 320422 17332
rect 554774 17320 554780 17332
rect 320416 17292 554780 17320
rect 320416 17280 320422 17292
rect 554774 17280 554780 17292
rect 554832 17280 554838 17332
rect 321646 17212 321652 17264
rect 321704 17252 321710 17264
rect 557534 17252 557540 17264
rect 321704 17224 557540 17252
rect 321704 17212 321710 17224
rect 557534 17212 557540 17224
rect 557592 17212 557598 17264
rect 241606 17144 241612 17196
rect 241664 17184 241670 17196
rect 362954 17184 362960 17196
rect 241664 17156 362960 17184
rect 241664 17144 241670 17156
rect 362954 17144 362960 17156
rect 363012 17144 363018 17196
rect 240226 17076 240232 17128
rect 240284 17116 240290 17128
rect 358814 17116 358820 17128
rect 240284 17088 358820 17116
rect 240284 17076 240290 17088
rect 358814 17076 358820 17088
rect 358872 17076 358878 17128
rect 237466 17008 237472 17060
rect 237524 17048 237530 17060
rect 356054 17048 356060 17060
rect 237524 17020 356060 17048
rect 237524 17008 237530 17020
rect 356054 17008 356060 17020
rect 356112 17008 356118 17060
rect 233418 16532 233424 16584
rect 233476 16572 233482 16584
rect 344554 16572 344560 16584
rect 233476 16544 344560 16572
rect 233476 16532 233482 16544
rect 344554 16532 344560 16544
rect 344612 16532 344618 16584
rect 313366 16464 313372 16516
rect 313424 16504 313430 16516
rect 539594 16504 539600 16516
rect 313424 16476 539600 16504
rect 313424 16464 313430 16476
rect 539594 16464 539600 16476
rect 539652 16464 539658 16516
rect 314838 16396 314844 16448
rect 314896 16436 314902 16448
rect 542722 16436 542728 16448
rect 314896 16408 542728 16436
rect 314896 16396 314902 16408
rect 542722 16396 542728 16408
rect 542780 16396 542786 16448
rect 316218 16328 316224 16380
rect 316276 16368 316282 16380
rect 546494 16368 546500 16380
rect 316276 16340 546500 16368
rect 316276 16328 316282 16340
rect 546494 16328 546500 16340
rect 546552 16328 546558 16380
rect 317506 16260 317512 16312
rect 317564 16300 317570 16312
rect 550266 16300 550272 16312
rect 317564 16272 550272 16300
rect 317564 16260 317570 16272
rect 550266 16260 550272 16272
rect 550324 16260 550330 16312
rect 318886 16192 318892 16244
rect 318944 16232 318950 16244
rect 553762 16232 553768 16244
rect 318944 16204 553768 16232
rect 318944 16192 318950 16204
rect 553762 16192 553768 16204
rect 553820 16192 553826 16244
rect 323118 16124 323124 16176
rect 323176 16164 323182 16176
rect 560386 16164 560392 16176
rect 323176 16136 560392 16164
rect 323176 16124 323182 16136
rect 560386 16124 560392 16136
rect 560444 16124 560450 16176
rect 324498 16056 324504 16108
rect 324556 16096 324562 16108
rect 564434 16096 564440 16108
rect 324556 16068 564440 16096
rect 324556 16056 324562 16068
rect 564434 16056 564440 16068
rect 564492 16056 564498 16108
rect 325786 15988 325792 16040
rect 325844 16028 325850 16040
rect 567562 16028 567568 16040
rect 325844 16000 567568 16028
rect 325844 15988 325850 16000
rect 567562 15988 567568 16000
rect 567620 15988 567626 16040
rect 327166 15920 327172 15972
rect 327224 15960 327230 15972
rect 571334 15960 571340 15972
rect 327224 15932 571340 15960
rect 327224 15920 327230 15932
rect 571334 15920 571340 15932
rect 571392 15920 571398 15972
rect 216858 15852 216864 15904
rect 216916 15892 216922 15904
rect 303890 15892 303896 15904
rect 216916 15864 303896 15892
rect 216916 15852 216922 15864
rect 303890 15852 303896 15864
rect 303948 15852 303954 15904
rect 328546 15852 328552 15904
rect 328604 15892 328610 15904
rect 575106 15892 575112 15904
rect 328604 15864 575112 15892
rect 328604 15852 328610 15864
rect 575106 15852 575112 15864
rect 575164 15852 575170 15904
rect 231946 15784 231952 15836
rect 232004 15824 232010 15836
rect 340966 15824 340972 15836
rect 232004 15796 340972 15824
rect 232004 15784 232010 15796
rect 340966 15784 340972 15796
rect 341024 15784 341030 15836
rect 230566 15716 230572 15768
rect 230624 15756 230630 15768
rect 337010 15756 337016 15768
rect 230624 15728 337016 15756
rect 230624 15716 230630 15728
rect 337010 15716 337016 15728
rect 337068 15716 337074 15768
rect 229186 15648 229192 15700
rect 229244 15688 229250 15700
rect 332686 15688 332692 15700
rect 229244 15660 332692 15688
rect 229244 15648 229250 15660
rect 332686 15648 332692 15660
rect 332744 15648 332750 15700
rect 289906 15104 289912 15156
rect 289964 15144 289970 15156
rect 482370 15144 482376 15156
rect 289964 15116 482376 15144
rect 289964 15104 289970 15116
rect 482370 15104 482376 15116
rect 482428 15104 482434 15156
rect 291286 15036 291292 15088
rect 291344 15076 291350 15088
rect 486418 15076 486424 15088
rect 291344 15048 486424 15076
rect 291344 15036 291350 15048
rect 486418 15036 486424 15048
rect 486476 15036 486482 15088
rect 292666 14968 292672 15020
rect 292724 15008 292730 15020
rect 490006 15008 490012 15020
rect 292724 14980 490012 15008
rect 292724 14968 292730 14980
rect 490006 14968 490012 14980
rect 490064 14968 490070 15020
rect 294046 14900 294052 14952
rect 294104 14940 294110 14952
rect 493042 14940 493048 14952
rect 294104 14912 493048 14940
rect 294104 14900 294110 14912
rect 493042 14900 493048 14912
rect 493100 14900 493106 14952
rect 298186 14832 298192 14884
rect 298244 14872 298250 14884
rect 500586 14872 500592 14884
rect 298244 14844 500592 14872
rect 298244 14832 298250 14844
rect 500586 14832 500592 14844
rect 500644 14832 500650 14884
rect 295426 14764 295432 14816
rect 295484 14804 295490 14816
rect 497090 14804 497096 14816
rect 295484 14776 497096 14804
rect 295484 14764 295490 14776
rect 497090 14764 497096 14776
rect 497148 14764 497154 14816
rect 299566 14696 299572 14748
rect 299624 14736 299630 14748
rect 503714 14736 503720 14748
rect 299624 14708 503720 14736
rect 299624 14696 299630 14708
rect 503714 14696 503720 14708
rect 503772 14696 503778 14748
rect 300946 14628 300952 14680
rect 301004 14668 301010 14680
rect 507210 14668 507216 14680
rect 301004 14640 507216 14668
rect 301004 14628 301010 14640
rect 507210 14628 507216 14640
rect 507268 14628 507274 14680
rect 302326 14560 302332 14612
rect 302384 14600 302390 14612
rect 511258 14600 511264 14612
rect 302384 14572 511264 14600
rect 302384 14560 302390 14572
rect 511258 14560 511264 14572
rect 511316 14560 511322 14612
rect 303706 14492 303712 14544
rect 303764 14532 303770 14544
rect 514754 14532 514760 14544
rect 303764 14504 514760 14532
rect 303764 14492 303770 14504
rect 514754 14492 514760 14504
rect 514812 14492 514818 14544
rect 305086 14424 305092 14476
rect 305144 14464 305150 14476
rect 517882 14464 517888 14476
rect 305144 14436 517888 14464
rect 305144 14424 305150 14436
rect 517882 14424 517888 14436
rect 517940 14424 517946 14476
rect 288526 14356 288532 14408
rect 288584 14396 288590 14408
rect 478138 14396 478144 14408
rect 288584 14368 478144 14396
rect 288584 14356 288590 14368
rect 478138 14356 478144 14368
rect 478196 14356 478202 14408
rect 287238 14288 287244 14340
rect 287296 14328 287302 14340
rect 474090 14328 474096 14340
rect 287296 14300 474096 14328
rect 287296 14288 287302 14300
rect 474090 14288 474096 14300
rect 474148 14288 474154 14340
rect 227806 14220 227812 14272
rect 227864 14260 227870 14272
rect 330386 14260 330392 14272
rect 227864 14232 330392 14260
rect 227864 14220 227870 14232
rect 330386 14220 330392 14232
rect 330444 14220 330450 14272
rect 263594 13744 263600 13796
rect 263652 13784 263658 13796
rect 417418 13784 417424 13796
rect 263652 13756 417424 13784
rect 263652 13744 263658 13756
rect 417418 13744 417424 13756
rect 417476 13744 417482 13796
rect 265066 13676 265072 13728
rect 265124 13716 265130 13728
rect 420914 13716 420920 13728
rect 265124 13688 420920 13716
rect 265124 13676 265130 13688
rect 420914 13676 420920 13688
rect 420972 13676 420978 13728
rect 266354 13608 266360 13660
rect 266412 13648 266418 13660
rect 423766 13648 423772 13660
rect 266412 13620 423772 13648
rect 266412 13608 266418 13620
rect 423766 13608 423772 13620
rect 423824 13608 423830 13660
rect 267734 13540 267740 13592
rect 267792 13580 267798 13592
rect 428458 13580 428464 13592
rect 267792 13552 428464 13580
rect 267792 13540 267798 13552
rect 428458 13540 428464 13552
rect 428516 13540 428522 13592
rect 269114 13472 269120 13524
rect 269172 13512 269178 13524
rect 432046 13512 432052 13524
rect 269172 13484 432052 13512
rect 269172 13472 269178 13484
rect 432046 13472 432052 13484
rect 432104 13472 432110 13524
rect 270494 13404 270500 13456
rect 270552 13444 270558 13456
rect 435082 13444 435088 13456
rect 270552 13416 435088 13444
rect 270552 13404 270558 13416
rect 435082 13404 435088 13416
rect 435140 13404 435146 13456
rect 271874 13336 271880 13388
rect 271932 13376 271938 13388
rect 439130 13376 439136 13388
rect 271932 13348 439136 13376
rect 271932 13336 271938 13348
rect 439130 13336 439136 13348
rect 439188 13336 439194 13388
rect 273438 13268 273444 13320
rect 273496 13308 273502 13320
rect 442626 13308 442632 13320
rect 273496 13280 442632 13308
rect 273496 13268 273502 13280
rect 442626 13268 442632 13280
rect 442684 13268 442690 13320
rect 274818 13200 274824 13252
rect 274876 13240 274882 13252
rect 445754 13240 445760 13252
rect 274876 13212 445760 13240
rect 274876 13200 274882 13212
rect 445754 13200 445760 13212
rect 445812 13200 445818 13252
rect 276198 13132 276204 13184
rect 276256 13172 276262 13184
rect 448514 13172 448520 13184
rect 276256 13144 448520 13172
rect 276256 13132 276262 13144
rect 448514 13132 448520 13144
rect 448572 13132 448578 13184
rect 277578 13064 277584 13116
rect 277636 13104 277642 13116
rect 453298 13104 453304 13116
rect 277636 13076 453304 13104
rect 277636 13064 277642 13076
rect 453298 13064 453304 13076
rect 453356 13064 453362 13116
rect 262306 12996 262312 13048
rect 262364 13036 262370 13048
rect 414290 13036 414296 13048
rect 262364 13008 414296 13036
rect 262364 12996 262370 13008
rect 414290 12996 414296 13008
rect 414348 12996 414354 13048
rect 260926 12928 260932 12980
rect 260984 12968 260990 12980
rect 410794 12968 410800 12980
rect 260984 12940 410800 12968
rect 260984 12928 260990 12940
rect 410794 12928 410800 12940
rect 410852 12928 410858 12980
rect 259546 12860 259552 12912
rect 259604 12900 259610 12912
rect 407206 12900 407212 12912
rect 259604 12872 407212 12900
rect 259604 12860 259610 12872
rect 407206 12860 407212 12872
rect 407264 12860 407270 12912
rect 236086 12384 236092 12436
rect 236144 12424 236150 12436
rect 349154 12424 349160 12436
rect 236144 12396 349160 12424
rect 236144 12384 236150 12396
rect 349154 12384 349160 12396
rect 349212 12384 349218 12436
rect 237374 12316 237380 12368
rect 237432 12356 237438 12368
rect 353570 12356 353576 12368
rect 237432 12328 353576 12356
rect 237432 12316 237438 12328
rect 353570 12316 353576 12328
rect 353628 12316 353634 12368
rect 238754 12248 238760 12300
rect 238812 12288 238818 12300
rect 357526 12288 357532 12300
rect 238812 12260 357532 12288
rect 238812 12248 238818 12260
rect 357526 12248 357532 12260
rect 357584 12248 357590 12300
rect 240134 12180 240140 12232
rect 240192 12220 240198 12232
rect 361114 12220 361120 12232
rect 240192 12192 361120 12220
rect 240192 12180 240198 12192
rect 361114 12180 361120 12192
rect 361172 12180 361178 12232
rect 241514 12112 241520 12164
rect 241572 12152 241578 12164
rect 364610 12152 364616 12164
rect 241572 12124 364616 12152
rect 241572 12112 241578 12124
rect 364610 12112 364616 12124
rect 364668 12112 364674 12164
rect 242894 12044 242900 12096
rect 242952 12084 242958 12096
rect 367738 12084 367744 12096
rect 242952 12056 367744 12084
rect 242952 12044 242958 12056
rect 367738 12044 367744 12056
rect 367796 12044 367802 12096
rect 244274 11976 244280 12028
rect 244332 12016 244338 12028
rect 371234 12016 371240 12028
rect 244332 11988 371240 12016
rect 244332 11976 244338 11988
rect 371234 11976 371240 11988
rect 371292 11976 371298 12028
rect 245746 11908 245752 11960
rect 245804 11948 245810 11960
rect 373994 11948 374000 11960
rect 245804 11920 374000 11948
rect 245804 11908 245810 11920
rect 373994 11908 374000 11920
rect 374052 11908 374058 11960
rect 247126 11840 247132 11892
rect 247184 11880 247190 11892
rect 378410 11880 378416 11892
rect 247184 11852 378416 11880
rect 247184 11840 247190 11852
rect 378410 11840 378416 11852
rect 378468 11840 378474 11892
rect 248506 11772 248512 11824
rect 248564 11812 248570 11824
rect 382366 11812 382372 11824
rect 248564 11784 382372 11812
rect 248564 11772 248570 11784
rect 382366 11772 382372 11784
rect 382424 11772 382430 11824
rect 249886 11704 249892 11756
rect 249944 11744 249950 11756
rect 385954 11744 385960 11756
rect 249944 11716 385960 11744
rect 249944 11704 249950 11716
rect 385954 11704 385960 11716
rect 386012 11704 386018 11756
rect 110414 11636 110420 11688
rect 110472 11676 110478 11688
rect 110598 11676 110604 11688
rect 110472 11648 110604 11676
rect 110472 11636 110478 11648
rect 110598 11636 110604 11648
rect 110656 11636 110662 11688
rect 234706 11636 234712 11688
rect 234764 11676 234770 11688
rect 346946 11676 346952 11688
rect 234764 11648 346952 11676
rect 234764 11636 234770 11648
rect 346946 11636 346952 11648
rect 347004 11636 347010 11688
rect 233326 11568 233332 11620
rect 233384 11608 233390 11620
rect 342898 11608 342904 11620
rect 233384 11580 342904 11608
rect 233384 11568 233390 11580
rect 342898 11568 342904 11580
rect 342956 11568 342962 11620
rect 226518 11500 226524 11552
rect 226576 11540 226582 11552
rect 326338 11540 326344 11552
rect 226576 11512 326344 11540
rect 226576 11500 226582 11512
rect 326338 11500 326344 11512
rect 326396 11500 326402 11552
rect 284294 11432 284300 11484
rect 284352 11472 284358 11484
rect 284478 11472 284484 11484
rect 284352 11444 284484 11472
rect 284352 11432 284358 11444
rect 284478 11432 284484 11444
rect 284536 11432 284542 11484
rect 309226 10956 309232 11008
rect 309284 10996 309290 11008
rect 527818 10996 527824 11008
rect 309284 10968 527824 10996
rect 309284 10956 309290 10968
rect 527818 10956 527824 10968
rect 527876 10956 527882 11008
rect 214098 10888 214104 10940
rect 214156 10928 214162 10940
rect 298186 10928 298192 10940
rect 214156 10900 298192 10928
rect 214156 10888 214162 10900
rect 298186 10888 298192 10900
rect 298244 10888 298250 10940
rect 310606 10888 310612 10940
rect 310664 10928 310670 10940
rect 531406 10928 531412 10940
rect 310664 10900 531412 10928
rect 310664 10888 310670 10900
rect 531406 10888 531412 10900
rect 531464 10888 531470 10940
rect 215478 10820 215484 10872
rect 215536 10860 215542 10872
rect 301498 10860 301504 10872
rect 215536 10832 301504 10860
rect 215536 10820 215542 10832
rect 301498 10820 301504 10832
rect 301556 10820 301562 10872
rect 311986 10820 311992 10872
rect 312044 10860 312050 10872
rect 534442 10860 534448 10872
rect 312044 10832 534448 10860
rect 312044 10820 312050 10832
rect 534442 10820 534448 10832
rect 534500 10820 534506 10872
rect 216766 10752 216772 10804
rect 216824 10792 216830 10804
rect 305546 10792 305552 10804
rect 216824 10764 305552 10792
rect 216824 10752 216830 10764
rect 305546 10752 305552 10764
rect 305604 10752 305610 10804
rect 313274 10752 313280 10804
rect 313332 10792 313338 10804
rect 538214 10792 538220 10804
rect 313332 10764 538220 10792
rect 313332 10752 313338 10764
rect 538214 10752 538220 10764
rect 538272 10752 538278 10804
rect 218238 10684 218244 10736
rect 218296 10724 218302 10736
rect 307938 10724 307944 10736
rect 218296 10696 307944 10724
rect 218296 10684 218302 10696
rect 307938 10684 307944 10696
rect 307996 10684 308002 10736
rect 314746 10684 314752 10736
rect 314804 10724 314810 10736
rect 541986 10724 541992 10736
rect 314804 10696 541992 10724
rect 314804 10684 314810 10696
rect 541986 10684 541992 10696
rect 542044 10684 542050 10736
rect 218146 10616 218152 10668
rect 218204 10656 218210 10668
rect 309042 10656 309048 10668
rect 218204 10628 309048 10656
rect 218204 10616 218210 10628
rect 309042 10616 309048 10628
rect 309100 10616 309106 10668
rect 316126 10616 316132 10668
rect 316184 10656 316190 10668
rect 545482 10656 545488 10668
rect 316184 10628 545488 10656
rect 316184 10616 316190 10628
rect 545482 10616 545488 10628
rect 545540 10616 545546 10668
rect 219526 10548 219532 10600
rect 219584 10588 219590 10600
rect 311434 10588 311440 10600
rect 219584 10560 311440 10588
rect 219584 10548 219590 10560
rect 311434 10548 311440 10560
rect 311492 10548 311498 10600
rect 317414 10548 317420 10600
rect 317472 10588 317478 10600
rect 548610 10588 548616 10600
rect 317472 10560 548616 10588
rect 317472 10548 317478 10560
rect 548610 10548 548616 10560
rect 548668 10548 548674 10600
rect 219618 10480 219624 10532
rect 219676 10520 219682 10532
rect 312170 10520 312176 10532
rect 219676 10492 312176 10520
rect 219676 10480 219682 10492
rect 312170 10480 312176 10492
rect 312228 10480 312234 10532
rect 318794 10480 318800 10532
rect 318852 10520 318858 10532
rect 552658 10520 552664 10532
rect 318852 10492 552664 10520
rect 318852 10480 318858 10492
rect 552658 10480 552664 10492
rect 552716 10480 552722 10532
rect 220998 10412 221004 10464
rect 221056 10452 221062 10464
rect 314746 10452 314752 10464
rect 221056 10424 314752 10452
rect 221056 10412 221062 10424
rect 314746 10412 314752 10424
rect 314804 10412 314810 10464
rect 320174 10412 320180 10464
rect 320232 10452 320238 10464
rect 556246 10452 556252 10464
rect 320232 10424 556252 10452
rect 320232 10412 320238 10424
rect 556246 10412 556252 10424
rect 556304 10412 556310 10464
rect 222194 10344 222200 10396
rect 222252 10384 222258 10396
rect 318058 10384 318064 10396
rect 222252 10356 318064 10384
rect 222252 10344 222258 10356
rect 318058 10344 318064 10356
rect 318116 10344 318122 10396
rect 323026 10344 323032 10396
rect 323084 10384 323090 10396
rect 563054 10384 563060 10396
rect 323084 10356 563060 10384
rect 323084 10344 323090 10356
rect 563054 10344 563060 10356
rect 563112 10344 563118 10396
rect 220906 10276 220912 10328
rect 220964 10316 220970 10328
rect 316218 10316 316224 10328
rect 220964 10288 316224 10316
rect 220964 10276 220970 10288
rect 316218 10276 316224 10288
rect 316276 10276 316282 10328
rect 324406 10276 324412 10328
rect 324464 10316 324470 10328
rect 566826 10316 566832 10328
rect 324464 10288 566832 10316
rect 324464 10276 324470 10288
rect 566826 10276 566832 10288
rect 566884 10276 566890 10328
rect 307846 10208 307852 10260
rect 307904 10248 307910 10260
rect 523770 10248 523776 10260
rect 307904 10220 523776 10248
rect 307904 10208 307910 10220
rect 523770 10208 523776 10220
rect 523828 10208 523834 10260
rect 306466 10140 306472 10192
rect 306524 10180 306530 10192
rect 520274 10180 520280 10192
rect 306524 10152 520280 10180
rect 306524 10140 306530 10152
rect 520274 10140 520280 10152
rect 520332 10140 520338 10192
rect 226426 10072 226432 10124
rect 226484 10112 226490 10124
rect 328730 10112 328736 10124
rect 226484 10084 328736 10112
rect 226484 10072 226490 10084
rect 328730 10072 328736 10084
rect 328788 10072 328794 10124
rect 225138 10004 225144 10056
rect 225196 10044 225202 10056
rect 324406 10044 324412 10056
rect 225196 10016 324412 10044
rect 225196 10004 225202 10016
rect 324406 10004 324412 10016
rect 324464 10004 324470 10056
rect 225046 9936 225052 9988
rect 225104 9976 225110 9988
rect 323026 9976 323032 9988
rect 225104 9948 323032 9976
rect 225104 9936 225110 9948
rect 323026 9936 323032 9948
rect 323084 9936 323090 9988
rect 223574 9868 223580 9920
rect 223632 9908 223638 9920
rect 319714 9908 319720 9920
rect 223632 9880 319720 9908
rect 223632 9868 223638 9880
rect 319714 9868 319720 9880
rect 319772 9868 319778 9920
rect 278866 9596 278872 9648
rect 278924 9636 278930 9648
rect 455690 9636 455696 9648
rect 278924 9608 455696 9636
rect 278924 9596 278930 9608
rect 455690 9596 455696 9608
rect 455748 9596 455754 9648
rect 280246 9528 280252 9580
rect 280304 9568 280310 9580
rect 459186 9568 459192 9580
rect 280304 9540 459192 9568
rect 280304 9528 280310 9540
rect 459186 9528 459192 9540
rect 459244 9528 459250 9580
rect 281626 9460 281632 9512
rect 281684 9500 281690 9512
rect 462774 9500 462780 9512
rect 281684 9472 462780 9500
rect 281684 9460 281690 9472
rect 462774 9460 462780 9472
rect 462832 9460 462838 9512
rect 283006 9392 283012 9444
rect 283064 9432 283070 9444
rect 466270 9432 466276 9444
rect 283064 9404 466276 9432
rect 283064 9392 283070 9404
rect 466270 9392 466276 9404
rect 466328 9392 466334 9444
rect 85666 9324 85672 9376
rect 85724 9364 85730 9376
rect 127158 9364 127164 9376
rect 85724 9336 127164 9364
rect 85724 9324 85730 9336
rect 127158 9324 127164 9336
rect 127216 9324 127222 9376
rect 203150 9324 203156 9376
rect 203208 9364 203214 9376
rect 270034 9364 270040 9376
rect 203208 9336 270040 9364
rect 203208 9324 203214 9336
rect 270034 9324 270040 9336
rect 270092 9324 270098 9376
rect 285766 9324 285772 9376
rect 285824 9364 285830 9376
rect 473446 9364 473452 9376
rect 285824 9336 473452 9364
rect 285824 9324 285830 9336
rect 473446 9324 473452 9336
rect 473504 9324 473510 9376
rect 45462 9256 45468 9308
rect 45520 9296 45526 9308
rect 110874 9296 110880 9308
rect 45520 9268 110880 9296
rect 45520 9256 45526 9268
rect 110874 9256 110880 9268
rect 110932 9256 110938 9308
rect 204254 9256 204260 9308
rect 204312 9296 204318 9308
rect 273622 9296 273628 9308
rect 204312 9268 273628 9296
rect 204312 9256 204318 9268
rect 273622 9256 273628 9268
rect 273680 9256 273686 9308
rect 287146 9256 287152 9308
rect 287204 9296 287210 9308
rect 476942 9296 476948 9308
rect 287204 9268 476948 9296
rect 287204 9256 287210 9268
rect 476942 9256 476948 9268
rect 477000 9256 477006 9308
rect 41874 9188 41880 9240
rect 41932 9228 41938 9240
rect 109126 9228 109132 9240
rect 41932 9200 109132 9228
rect 41932 9188 41938 9200
rect 109126 9188 109132 9200
rect 109184 9188 109190 9240
rect 205634 9188 205640 9240
rect 205692 9228 205698 9240
rect 277118 9228 277124 9240
rect 205692 9200 277124 9228
rect 205692 9188 205698 9200
rect 277118 9188 277124 9200
rect 277176 9188 277182 9240
rect 289814 9188 289820 9240
rect 289872 9228 289878 9240
rect 481726 9228 481732 9240
rect 289872 9200 481732 9228
rect 289872 9188 289878 9200
rect 481726 9188 481732 9200
rect 481784 9188 481790 9240
rect 38378 9120 38384 9172
rect 38436 9160 38442 9172
rect 107838 9160 107844 9172
rect 38436 9132 107844 9160
rect 38436 9120 38442 9132
rect 107838 9120 107844 9132
rect 107896 9120 107902 9172
rect 207106 9120 207112 9172
rect 207164 9160 207170 9172
rect 280706 9160 280712 9172
rect 207164 9132 280712 9160
rect 207164 9120 207170 9132
rect 280706 9120 280712 9132
rect 280764 9120 280770 9172
rect 291194 9120 291200 9172
rect 291252 9160 291258 9172
rect 485222 9160 485228 9172
rect 291252 9132 485228 9160
rect 291252 9120 291258 9132
rect 485222 9120 485228 9132
rect 485280 9120 485286 9172
rect 34790 9052 34796 9104
rect 34848 9092 34854 9104
rect 106458 9092 106464 9104
rect 34848 9064 106464 9092
rect 34848 9052 34854 9064
rect 106458 9052 106464 9064
rect 106516 9052 106522 9104
rect 208486 9052 208492 9104
rect 208544 9092 208550 9104
rect 284294 9092 284300 9104
rect 208544 9064 284300 9092
rect 208544 9052 208550 9064
rect 284294 9052 284300 9064
rect 284352 9052 284358 9104
rect 292574 9052 292580 9104
rect 292632 9092 292638 9104
rect 488810 9092 488816 9104
rect 292632 9064 488816 9092
rect 292632 9052 292638 9064
rect 488810 9052 488816 9064
rect 488868 9052 488874 9104
rect 31294 8984 31300 9036
rect 31352 9024 31358 9036
rect 103606 9024 103612 9036
rect 31352 8996 103612 9024
rect 31352 8984 31358 8996
rect 103606 8984 103612 8996
rect 103664 8984 103670 9036
rect 209866 8984 209872 9036
rect 209924 9024 209930 9036
rect 287790 9024 287796 9036
rect 209924 8996 287796 9024
rect 209924 8984 209930 8996
rect 287790 8984 287796 8996
rect 287848 8984 287854 9036
rect 293954 8984 293960 9036
rect 294012 9024 294018 9036
rect 492306 9024 492312 9036
rect 294012 8996 492312 9024
rect 294012 8984 294018 8996
rect 492306 8984 492312 8996
rect 492364 8984 492370 9036
rect 27706 8916 27712 8968
rect 27764 8956 27770 8968
rect 102226 8956 102232 8968
rect 27764 8928 102232 8956
rect 27764 8916 27770 8928
rect 102226 8916 102232 8928
rect 102284 8916 102290 8968
rect 211246 8916 211252 8968
rect 211304 8956 211310 8968
rect 291378 8956 291384 8968
rect 211304 8928 291384 8956
rect 211304 8916 211310 8928
rect 291378 8916 291384 8928
rect 291436 8916 291442 8968
rect 296806 8916 296812 8968
rect 296864 8956 296870 8968
rect 499390 8956 499396 8968
rect 296864 8928 499396 8956
rect 296864 8916 296870 8928
rect 499390 8916 499396 8928
rect 499448 8916 499454 8968
rect 276106 8848 276112 8900
rect 276164 8888 276170 8900
rect 448606 8888 448612 8900
rect 276164 8860 448612 8888
rect 276164 8848 276170 8860
rect 448606 8848 448612 8860
rect 448664 8848 448670 8900
rect 273346 8780 273352 8832
rect 273404 8820 273410 8832
rect 441522 8820 441528 8832
rect 273404 8792 441528 8820
rect 273404 8780 273410 8792
rect 441522 8780 441528 8792
rect 441580 8780 441586 8832
rect 215386 8712 215392 8764
rect 215444 8752 215450 8764
rect 300762 8752 300768 8764
rect 215444 8724 300768 8752
rect 215444 8712 215450 8724
rect 300762 8712 300768 8724
rect 300820 8712 300826 8764
rect 214006 8644 214012 8696
rect 214064 8684 214070 8696
rect 297266 8684 297272 8696
rect 214064 8656 297272 8684
rect 214064 8644 214070 8656
rect 297266 8644 297272 8656
rect 297324 8644 297330 8696
rect 212534 8576 212540 8628
rect 212592 8616 212598 8628
rect 294874 8616 294880 8628
rect 212592 8588 294880 8616
rect 212592 8576 212598 8588
rect 294874 8576 294880 8588
rect 294932 8576 294938 8628
rect 51350 8236 51356 8288
rect 51408 8276 51414 8288
rect 111978 8276 111984 8288
rect 51408 8248 111984 8276
rect 51408 8236 51414 8248
rect 111978 8236 111984 8248
rect 112036 8236 112042 8288
rect 249794 8236 249800 8288
rect 249852 8276 249858 8288
rect 384758 8276 384764 8288
rect 249852 8248 384764 8276
rect 249852 8236 249858 8248
rect 384758 8236 384764 8248
rect 384816 8236 384822 8288
rect 47854 8168 47860 8220
rect 47912 8208 47918 8220
rect 110782 8208 110788 8220
rect 47912 8180 110788 8208
rect 47912 8168 47918 8180
rect 110782 8168 110788 8180
rect 110840 8168 110846 8220
rect 251174 8168 251180 8220
rect 251232 8208 251238 8220
rect 388254 8208 388260 8220
rect 251232 8180 388260 8208
rect 251232 8168 251238 8180
rect 388254 8168 388260 8180
rect 388312 8168 388318 8220
rect 33594 8100 33600 8152
rect 33652 8140 33658 8152
rect 105078 8140 105084 8152
rect 33652 8112 105084 8140
rect 33652 8100 33658 8112
rect 105078 8100 105084 8112
rect 105136 8100 105142 8152
rect 201586 8100 201592 8152
rect 201644 8140 201650 8152
rect 237374 8140 237380 8152
rect 201644 8112 237380 8140
rect 201644 8100 201650 8112
rect 237374 8100 237380 8112
rect 237432 8100 237438 8152
rect 252554 8100 252560 8152
rect 252612 8140 252618 8152
rect 391842 8140 391848 8152
rect 252612 8112 391848 8140
rect 252612 8100 252618 8112
rect 391842 8100 391848 8112
rect 391900 8100 391906 8152
rect 30098 8032 30104 8084
rect 30156 8072 30162 8084
rect 103698 8072 103704 8084
rect 30156 8044 103704 8072
rect 30156 8032 30162 8044
rect 103698 8032 103704 8044
rect 103756 8032 103762 8084
rect 203058 8032 203064 8084
rect 203116 8072 203122 8084
rect 240134 8072 240140 8084
rect 203116 8044 240140 8072
rect 203116 8032 203122 8044
rect 240134 8032 240140 8044
rect 240192 8032 240198 8084
rect 253934 8032 253940 8084
rect 253992 8072 253998 8084
rect 395338 8072 395344 8084
rect 253992 8044 395344 8072
rect 253992 8032 253998 8044
rect 395338 8032 395344 8044
rect 395396 8032 395402 8084
rect 26510 7964 26516 8016
rect 26568 8004 26574 8016
rect 102318 8004 102324 8016
rect 26568 7976 102324 8004
rect 26568 7964 26574 7976
rect 102318 7964 102324 7976
rect 102376 7964 102382 8016
rect 207014 7964 207020 8016
rect 207072 8004 207078 8016
rect 249794 8004 249800 8016
rect 207072 7976 249800 8004
rect 207072 7964 207078 7976
rect 249794 7964 249800 7976
rect 249852 7964 249858 8016
rect 255314 7964 255320 8016
rect 255372 8004 255378 8016
rect 398926 8004 398932 8016
rect 255372 7976 398932 8004
rect 255372 7964 255378 7976
rect 398926 7964 398932 7976
rect 398984 7964 398990 8016
rect 23014 7896 23020 7948
rect 23072 7936 23078 7948
rect 100938 7936 100944 7948
rect 23072 7908 100944 7936
rect 23072 7896 23078 7908
rect 100938 7896 100944 7908
rect 100996 7896 101002 7948
rect 187786 7896 187792 7948
rect 187844 7936 187850 7948
rect 234706 7936 234712 7948
rect 187844 7908 234712 7936
rect 187844 7896 187850 7908
rect 234706 7896 234712 7908
rect 234764 7896 234770 7948
rect 256694 7896 256700 7948
rect 256752 7936 256758 7948
rect 402514 7936 402520 7948
rect 256752 7908 402520 7936
rect 256752 7896 256758 7908
rect 402514 7896 402520 7908
rect 402572 7896 402578 7948
rect 18230 7828 18236 7880
rect 18288 7868 18294 7880
rect 99466 7868 99472 7880
rect 18288 7840 99472 7868
rect 18288 7828 18294 7840
rect 99466 7828 99472 7840
rect 99524 7828 99530 7880
rect 193490 7828 193496 7880
rect 193548 7868 193554 7880
rect 248782 7868 248788 7880
rect 193548 7840 248788 7868
rect 193548 7828 193554 7840
rect 248782 7828 248788 7840
rect 248840 7828 248846 7880
rect 258074 7828 258080 7880
rect 258132 7868 258138 7880
rect 406010 7868 406016 7880
rect 258132 7840 406016 7868
rect 258132 7828 258138 7840
rect 406010 7828 406016 7840
rect 406068 7828 406074 7880
rect 7650 7760 7656 7812
rect 7708 7800 7714 7812
rect 94038 7800 94044 7812
rect 7708 7772 94044 7800
rect 7708 7760 7714 7772
rect 94038 7760 94044 7772
rect 94096 7760 94102 7812
rect 194686 7760 194692 7812
rect 194744 7800 194750 7812
rect 251174 7800 251180 7812
rect 194744 7772 251180 7800
rect 194744 7760 194750 7772
rect 251174 7760 251180 7772
rect 251232 7760 251238 7812
rect 259454 7760 259460 7812
rect 259512 7800 259518 7812
rect 409598 7800 409604 7812
rect 259512 7772 409604 7800
rect 259512 7760 259518 7772
rect 409598 7760 409604 7772
rect 409656 7760 409662 7812
rect 2866 7692 2872 7744
rect 2924 7732 2930 7744
rect 92658 7732 92664 7744
rect 2924 7704 92664 7732
rect 2924 7692 2930 7704
rect 92658 7692 92664 7704
rect 92716 7692 92722 7744
rect 201494 7692 201500 7744
rect 201552 7732 201558 7744
rect 258074 7732 258080 7744
rect 201552 7704 258080 7732
rect 201552 7692 201558 7704
rect 258074 7692 258080 7704
rect 258132 7692 258138 7744
rect 260834 7692 260840 7744
rect 260892 7732 260898 7744
rect 413094 7732 413100 7744
rect 260892 7704 413100 7732
rect 260892 7692 260898 7704
rect 413094 7692 413100 7704
rect 413152 7692 413158 7744
rect 566 7624 572 7676
rect 624 7664 630 7676
rect 91094 7664 91100 7676
rect 624 7636 91100 7664
rect 624 7624 630 7636
rect 91094 7624 91100 7636
rect 91152 7624 91158 7676
rect 91554 7624 91560 7676
rect 91612 7664 91618 7676
rect 128538 7664 128544 7676
rect 91612 7636 128544 7664
rect 91612 7624 91618 7636
rect 128538 7624 128544 7636
rect 128596 7624 128602 7676
rect 197538 7624 197544 7676
rect 197596 7664 197602 7676
rect 255866 7664 255872 7676
rect 197596 7636 255872 7664
rect 197596 7624 197602 7636
rect 255866 7624 255872 7636
rect 255924 7624 255930 7676
rect 262214 7624 262220 7676
rect 262272 7664 262278 7676
rect 416682 7664 416688 7676
rect 262272 7636 416688 7664
rect 262272 7624 262278 7636
rect 416682 7624 416688 7636
rect 416740 7624 416746 7676
rect 1670 7556 1676 7608
rect 1728 7596 1734 7608
rect 92750 7596 92756 7608
rect 1728 7568 92756 7596
rect 1728 7556 1734 7568
rect 92750 7556 92756 7568
rect 92808 7556 92814 7608
rect 98638 7556 98644 7608
rect 98696 7596 98702 7608
rect 132586 7596 132592 7608
rect 98696 7568 132592 7596
rect 98696 7556 98702 7568
rect 132586 7556 132592 7568
rect 132644 7556 132650 7608
rect 198918 7556 198924 7608
rect 198976 7596 198982 7608
rect 261754 7596 261760 7608
rect 198976 7568 261760 7596
rect 198976 7556 198982 7568
rect 261754 7556 261760 7568
rect 261812 7556 261818 7608
rect 264974 7556 264980 7608
rect 265032 7596 265038 7608
rect 420178 7596 420184 7608
rect 265032 7568 420184 7596
rect 265032 7556 265038 7568
rect 420178 7556 420184 7568
rect 420236 7556 420242 7608
rect 54938 7488 54944 7540
rect 54996 7528 55002 7540
rect 114646 7528 114652 7540
rect 54996 7500 114652 7528
rect 54996 7488 55002 7500
rect 114646 7488 114652 7500
rect 114704 7488 114710 7540
rect 248414 7488 248420 7540
rect 248472 7528 248478 7540
rect 381170 7528 381176 7540
rect 248472 7500 381176 7528
rect 248472 7488 248478 7500
rect 381170 7488 381176 7500
rect 381228 7488 381234 7540
rect 84470 7420 84476 7472
rect 84528 7460 84534 7472
rect 125778 7460 125784 7472
rect 84528 7432 125784 7460
rect 84528 7420 84534 7432
rect 125778 7420 125784 7432
rect 125836 7420 125842 7472
rect 247034 7420 247040 7472
rect 247092 7460 247098 7472
rect 377674 7460 377680 7472
rect 247092 7432 377680 7460
rect 247092 7420 247098 7432
rect 377674 7420 377680 7432
rect 377732 7420 377738 7472
rect 87966 7352 87972 7404
rect 88024 7392 88030 7404
rect 127066 7392 127072 7404
rect 88024 7364 127072 7392
rect 88024 7352 88030 7364
rect 127066 7352 127072 7364
rect 127124 7352 127130 7404
rect 245654 7352 245660 7404
rect 245712 7392 245718 7404
rect 374086 7392 374092 7404
rect 245712 7364 374092 7392
rect 245712 7352 245718 7364
rect 374086 7352 374092 7364
rect 374144 7352 374150 7404
rect 200206 7284 200212 7336
rect 200264 7324 200270 7336
rect 265342 7324 265348 7336
rect 200264 7296 265348 7324
rect 200264 7284 200270 7296
rect 265342 7284 265348 7296
rect 265400 7284 265406 7336
rect 200298 7216 200304 7268
rect 200356 7256 200362 7268
rect 262950 7256 262956 7268
rect 200356 7228 262956 7256
rect 200356 7216 200362 7228
rect 262950 7216 262956 7228
rect 263008 7216 263014 7268
rect 73798 6808 73804 6860
rect 73856 6848 73862 6860
rect 121638 6848 121644 6860
rect 73856 6820 121644 6848
rect 73856 6808 73862 6820
rect 121638 6808 121644 6820
rect 121696 6808 121702 6860
rect 185026 6808 185032 6860
rect 185084 6848 185090 6860
rect 227530 6848 227536 6860
rect 185084 6820 227536 6848
rect 185084 6808 185090 6820
rect 227530 6808 227536 6820
rect 227588 6808 227594 6860
rect 231854 6808 231860 6860
rect 231912 6848 231918 6860
rect 342162 6848 342168 6860
rect 231912 6820 342168 6848
rect 231912 6808 231918 6820
rect 342162 6808 342168 6820
rect 342220 6808 342226 6860
rect 70302 6740 70308 6792
rect 70360 6780 70366 6792
rect 120166 6780 120172 6792
rect 70360 6752 120172 6780
rect 70360 6740 70366 6752
rect 120166 6740 120172 6752
rect 120224 6740 120230 6792
rect 185118 6740 185124 6792
rect 185176 6780 185182 6792
rect 226426 6780 226432 6792
rect 185176 6752 226432 6780
rect 185176 6740 185182 6752
rect 226426 6740 226432 6752
rect 226484 6740 226490 6792
rect 233234 6740 233240 6792
rect 233292 6780 233298 6792
rect 345750 6780 345756 6792
rect 233292 6752 345756 6780
rect 233292 6740 233298 6752
rect 345750 6740 345756 6752
rect 345808 6740 345814 6792
rect 66714 6672 66720 6724
rect 66772 6712 66778 6724
rect 118878 6712 118884 6724
rect 66772 6684 118884 6712
rect 66772 6672 66778 6684
rect 118878 6672 118884 6684
rect 118936 6672 118942 6724
rect 186498 6672 186504 6724
rect 186556 6712 186562 6724
rect 229830 6712 229836 6724
rect 186556 6684 229836 6712
rect 186556 6672 186562 6684
rect 229830 6672 229836 6684
rect 229888 6672 229894 6724
rect 234614 6672 234620 6724
rect 234672 6712 234678 6724
rect 349246 6712 349252 6724
rect 234672 6684 349252 6712
rect 234672 6672 234678 6684
rect 349246 6672 349252 6684
rect 349304 6672 349310 6724
rect 63218 6604 63224 6656
rect 63276 6644 63282 6656
rect 117498 6644 117504 6656
rect 63276 6616 117504 6644
rect 63276 6604 63282 6616
rect 117498 6604 117504 6616
rect 117556 6604 117562 6656
rect 187694 6604 187700 6656
rect 187752 6644 187758 6656
rect 233418 6644 233424 6656
rect 187752 6616 233424 6644
rect 187752 6604 187758 6616
rect 233418 6604 233424 6616
rect 233476 6604 233482 6656
rect 274726 6604 274732 6656
rect 274784 6644 274790 6656
rect 445018 6644 445024 6656
rect 274784 6616 445024 6644
rect 274784 6604 274790 6616
rect 445018 6604 445024 6616
rect 445076 6604 445082 6656
rect 59630 6536 59636 6588
rect 59688 6576 59694 6588
rect 116210 6576 116216 6588
rect 59688 6548 116216 6576
rect 59688 6536 59694 6548
rect 116210 6536 116216 6548
rect 116268 6536 116274 6588
rect 189350 6536 189356 6588
rect 189408 6576 189414 6588
rect 237006 6576 237012 6588
rect 189408 6548 237012 6576
rect 189408 6536 189414 6548
rect 237006 6536 237012 6548
rect 237064 6536 237070 6588
rect 277486 6536 277492 6588
rect 277544 6576 277550 6588
rect 452102 6576 452108 6588
rect 277544 6548 452108 6576
rect 277544 6536 277550 6548
rect 452102 6536 452108 6548
rect 452160 6536 452166 6588
rect 56042 6468 56048 6520
rect 56100 6508 56106 6520
rect 114738 6508 114744 6520
rect 56100 6480 114744 6508
rect 56100 6468 56106 6480
rect 114738 6468 114744 6480
rect 114796 6468 114802 6520
rect 190638 6468 190644 6520
rect 190696 6508 190702 6520
rect 240502 6508 240508 6520
rect 190696 6480 240508 6508
rect 190696 6468 190702 6480
rect 240502 6468 240508 6480
rect 240560 6468 240566 6520
rect 284386 6468 284392 6520
rect 284444 6508 284450 6520
rect 469858 6508 469864 6520
rect 284444 6480 469864 6508
rect 284444 6468 284450 6480
rect 469858 6468 469864 6480
rect 469916 6468 469922 6520
rect 52546 6400 52552 6452
rect 52604 6440 52610 6452
rect 113266 6440 113272 6452
rect 52604 6412 113272 6440
rect 52604 6400 52610 6412
rect 113266 6400 113272 6412
rect 113324 6400 113330 6452
rect 193398 6400 193404 6452
rect 193456 6440 193462 6452
rect 247586 6440 247592 6452
rect 193456 6412 247592 6440
rect 193456 6400 193462 6412
rect 247586 6400 247592 6412
rect 247644 6400 247650 6452
rect 322934 6400 322940 6452
rect 322992 6440 322998 6452
rect 562042 6440 562048 6452
rect 322992 6412 562048 6440
rect 322992 6400 322998 6412
rect 562042 6400 562048 6412
rect 562100 6400 562106 6452
rect 48958 6332 48964 6384
rect 49016 6372 49022 6384
rect 111886 6372 111892 6384
rect 49016 6344 111892 6372
rect 49016 6332 49022 6344
rect 111886 6332 111892 6344
rect 111944 6332 111950 6384
rect 196066 6332 196072 6384
rect 196124 6372 196130 6384
rect 254670 6372 254676 6384
rect 196124 6344 254676 6372
rect 196124 6332 196130 6344
rect 254670 6332 254676 6344
rect 254728 6332 254734 6384
rect 324314 6332 324320 6384
rect 324372 6372 324378 6384
rect 565630 6372 565636 6384
rect 324372 6344 565636 6372
rect 324372 6332 324378 6344
rect 565630 6332 565636 6344
rect 565688 6332 565694 6384
rect 44266 6264 44272 6316
rect 44324 6304 44330 6316
rect 109218 6304 109224 6316
rect 44324 6276 109224 6304
rect 44324 6264 44330 6276
rect 109218 6264 109224 6276
rect 109276 6264 109282 6316
rect 197446 6264 197452 6316
rect 197504 6304 197510 6316
rect 258258 6304 258264 6316
rect 197504 6276 258264 6304
rect 197504 6264 197510 6276
rect 258258 6264 258264 6276
rect 258316 6264 258322 6316
rect 325694 6264 325700 6316
rect 325752 6304 325758 6316
rect 569126 6304 569132 6316
rect 325752 6276 569132 6304
rect 325752 6264 325758 6276
rect 569126 6264 569132 6276
rect 569184 6264 569190 6316
rect 40678 6196 40684 6248
rect 40736 6236 40742 6248
rect 107746 6236 107752 6248
rect 40736 6208 107752 6236
rect 40736 6196 40742 6208
rect 107746 6196 107752 6208
rect 107804 6196 107810 6248
rect 192018 6196 192024 6248
rect 192076 6236 192082 6248
rect 244090 6236 244096 6248
rect 192076 6208 244096 6236
rect 192076 6196 192082 6208
rect 244090 6196 244096 6208
rect 244148 6196 244154 6248
rect 246298 6196 246304 6248
rect 246356 6236 246362 6248
rect 322106 6236 322112 6248
rect 246356 6208 322112 6236
rect 246356 6196 246362 6208
rect 322106 6196 322112 6208
rect 322164 6196 322170 6248
rect 327074 6196 327080 6248
rect 327132 6236 327138 6248
rect 572714 6236 572720 6248
rect 327132 6208 572720 6236
rect 327132 6196 327138 6208
rect 572714 6196 572720 6208
rect 572772 6196 572778 6248
rect 37182 6128 37188 6180
rect 37240 6168 37246 6180
rect 106366 6168 106372 6180
rect 37240 6140 106372 6168
rect 37240 6128 37246 6140
rect 106366 6128 106372 6140
rect 106424 6128 106430 6180
rect 183830 6128 183836 6180
rect 183888 6168 183894 6180
rect 222746 6168 222752 6180
rect 183888 6140 222752 6168
rect 183888 6128 183894 6140
rect 222746 6128 222752 6140
rect 222804 6128 222810 6180
rect 224954 6128 224960 6180
rect 225012 6168 225018 6180
rect 324314 6168 324320 6180
rect 225012 6140 324320 6168
rect 225012 6128 225018 6140
rect 324314 6128 324320 6140
rect 324372 6128 324378 6180
rect 328454 6128 328460 6180
rect 328512 6168 328518 6180
rect 576302 6168 576308 6180
rect 328512 6140 576308 6168
rect 328512 6128 328518 6140
rect 576302 6128 576308 6140
rect 576360 6128 576366 6180
rect 77386 6060 77392 6112
rect 77444 6100 77450 6112
rect 123018 6100 123024 6112
rect 77444 6072 123024 6100
rect 77444 6060 77450 6072
rect 123018 6060 123024 6072
rect 123076 6060 123082 6112
rect 180886 6060 180892 6112
rect 180944 6100 180950 6112
rect 215662 6100 215668 6112
rect 180944 6072 215668 6100
rect 180944 6060 180950 6072
rect 215662 6060 215668 6072
rect 215720 6060 215726 6112
rect 230474 6060 230480 6112
rect 230532 6100 230538 6112
rect 338666 6100 338672 6112
rect 230532 6072 338672 6100
rect 230532 6060 230538 6072
rect 338666 6060 338672 6072
rect 338724 6060 338730 6112
rect 80882 5992 80888 6044
rect 80940 6032 80946 6044
rect 124398 6032 124404 6044
rect 80940 6004 124404 6032
rect 80940 5992 80946 6004
rect 124398 5992 124404 6004
rect 124456 5992 124462 6044
rect 186406 5992 186412 6044
rect 186464 6032 186470 6044
rect 218054 6032 218060 6044
rect 186464 6004 218060 6032
rect 186464 5992 186470 6004
rect 218054 5992 218060 6004
rect 218112 5992 218118 6044
rect 229094 5992 229100 6044
rect 229152 6032 229158 6044
rect 335078 6032 335084 6044
rect 229152 6004 335084 6032
rect 229152 5992 229158 6004
rect 335078 5992 335084 6004
rect 335136 5992 335142 6044
rect 95142 5924 95148 5976
rect 95200 5964 95206 5976
rect 131298 5964 131304 5976
rect 95200 5936 131304 5964
rect 95200 5924 95206 5936
rect 131298 5924 131304 5936
rect 131356 5924 131362 5976
rect 185210 5924 185216 5976
rect 185268 5964 185274 5976
rect 216766 5964 216772 5976
rect 185268 5936 216772 5964
rect 185268 5924 185274 5936
rect 216766 5924 216772 5936
rect 216824 5924 216830 5976
rect 227714 5924 227720 5976
rect 227772 5964 227778 5976
rect 331582 5964 331588 5976
rect 227772 5936 331588 5964
rect 227772 5924 227778 5936
rect 331582 5924 331588 5936
rect 331640 5924 331646 5976
rect 333238 5924 333244 5976
rect 333296 5964 333302 5976
rect 418982 5964 418988 5976
rect 333296 5936 418988 5964
rect 333296 5924 333302 5936
rect 418982 5924 418988 5936
rect 419040 5924 419046 5976
rect 226334 5856 226340 5908
rect 226392 5896 226398 5908
rect 327994 5896 328000 5908
rect 226392 5868 328000 5896
rect 226392 5856 226398 5868
rect 327994 5856 328000 5868
rect 328052 5856 328058 5908
rect 243630 5788 243636 5840
rect 243688 5828 243694 5840
rect 293678 5828 293684 5840
rect 243688 5800 293684 5828
rect 243688 5788 243694 5800
rect 293678 5788 293684 5800
rect 293736 5788 293742 5840
rect 238018 5720 238024 5772
rect 238076 5760 238082 5772
rect 283098 5760 283104 5772
rect 238076 5732 283104 5760
rect 238076 5720 238082 5732
rect 283098 5720 283104 5732
rect 283156 5720 283162 5772
rect 79686 5448 79692 5500
rect 79744 5488 79750 5500
rect 124306 5488 124312 5500
rect 79744 5460 124312 5488
rect 79744 5448 79750 5460
rect 124306 5448 124312 5460
rect 124364 5448 124370 5500
rect 197354 5448 197360 5500
rect 197412 5488 197418 5500
rect 257062 5488 257068 5500
rect 197412 5460 257068 5488
rect 197412 5448 197418 5460
rect 257062 5448 257068 5460
rect 257120 5448 257126 5500
rect 257338 5448 257344 5500
rect 257396 5488 257402 5500
rect 290182 5488 290188 5500
rect 257396 5460 290188 5488
rect 257396 5448 257402 5460
rect 290182 5448 290188 5460
rect 290240 5448 290246 5500
rect 299474 5448 299480 5500
rect 299532 5488 299538 5500
rect 505370 5488 505376 5500
rect 299532 5460 505376 5488
rect 299532 5448 299538 5460
rect 505370 5448 505376 5460
rect 505428 5448 505434 5500
rect 76190 5380 76196 5432
rect 76248 5420 76254 5432
rect 122926 5420 122932 5432
rect 76248 5392 122932 5420
rect 76248 5380 76254 5392
rect 122926 5380 122932 5392
rect 122984 5380 122990 5432
rect 168466 5380 168472 5432
rect 168524 5420 168530 5432
rect 187326 5420 187332 5432
rect 168524 5392 187332 5420
rect 168524 5380 168530 5392
rect 187326 5380 187332 5392
rect 187384 5380 187390 5432
rect 198826 5380 198832 5432
rect 198884 5420 198890 5432
rect 260650 5420 260656 5432
rect 198884 5392 260656 5420
rect 198884 5380 198890 5392
rect 260650 5380 260656 5392
rect 260708 5380 260714 5432
rect 300854 5380 300860 5432
rect 300912 5420 300918 5432
rect 508866 5420 508872 5432
rect 300912 5392 508872 5420
rect 300912 5380 300918 5392
rect 508866 5380 508872 5392
rect 508924 5380 508930 5432
rect 72602 5312 72608 5364
rect 72660 5352 72666 5364
rect 121546 5352 121552 5364
rect 72660 5324 121552 5352
rect 72660 5312 72666 5324
rect 121546 5312 121552 5324
rect 121604 5312 121610 5364
rect 169938 5312 169944 5364
rect 169996 5352 170002 5364
rect 190822 5352 190828 5364
rect 169996 5324 190828 5352
rect 169996 5312 170002 5324
rect 190822 5312 190828 5324
rect 190880 5312 190886 5364
rect 202966 5312 202972 5364
rect 203024 5352 203030 5364
rect 271230 5352 271236 5364
rect 203024 5324 271236 5352
rect 203024 5312 203030 5324
rect 271230 5312 271236 5324
rect 271288 5312 271294 5364
rect 302234 5312 302240 5364
rect 302292 5352 302298 5364
rect 512454 5352 512460 5364
rect 302292 5324 512460 5352
rect 302292 5312 302298 5324
rect 512454 5312 512460 5324
rect 512512 5312 512518 5364
rect 69106 5244 69112 5296
rect 69164 5284 69170 5296
rect 120258 5284 120264 5296
rect 69164 5256 120264 5284
rect 69164 5244 69170 5256
rect 120258 5244 120264 5256
rect 120316 5244 120322 5296
rect 171134 5244 171140 5296
rect 171192 5284 171198 5296
rect 194410 5284 194416 5296
rect 171192 5256 194416 5284
rect 171192 5244 171198 5256
rect 194410 5244 194416 5256
rect 194468 5244 194474 5296
rect 208394 5244 208400 5296
rect 208452 5284 208458 5296
rect 285398 5284 285404 5296
rect 208452 5256 285404 5284
rect 208452 5244 208458 5256
rect 285398 5244 285404 5256
rect 285456 5244 285462 5296
rect 303614 5244 303620 5296
rect 303672 5284 303678 5296
rect 515950 5284 515956 5296
rect 303672 5256 515956 5284
rect 303672 5244 303678 5256
rect 515950 5244 515956 5256
rect 516008 5244 516014 5296
rect 62022 5176 62028 5228
rect 62080 5216 62086 5228
rect 117406 5216 117412 5228
rect 62080 5188 117412 5216
rect 62080 5176 62086 5188
rect 117406 5176 117412 5188
rect 117464 5176 117470 5228
rect 172606 5176 172612 5228
rect 172664 5216 172670 5228
rect 197906 5216 197912 5228
rect 172664 5188 197912 5216
rect 172664 5176 172670 5188
rect 197906 5176 197912 5188
rect 197964 5176 197970 5228
rect 209774 5176 209780 5228
rect 209832 5216 209838 5228
rect 288986 5216 288992 5228
rect 209832 5188 288992 5216
rect 209832 5176 209838 5188
rect 288986 5176 288992 5188
rect 289044 5176 289050 5228
rect 304994 5176 305000 5228
rect 305052 5216 305058 5228
rect 519538 5216 519544 5228
rect 305052 5188 519544 5216
rect 305052 5176 305058 5188
rect 519538 5176 519544 5188
rect 519596 5176 519602 5228
rect 58434 5108 58440 5160
rect 58492 5148 58498 5160
rect 116118 5148 116124 5160
rect 58492 5120 116124 5148
rect 58492 5108 58498 5120
rect 116118 5108 116124 5120
rect 116176 5108 116182 5160
rect 117222 5108 117228 5160
rect 117280 5148 117286 5160
rect 136818 5148 136824 5160
rect 117280 5120 136824 5148
rect 117280 5108 117286 5120
rect 136818 5108 136824 5120
rect 136876 5108 136882 5160
rect 173986 5108 173992 5160
rect 174044 5148 174050 5160
rect 201494 5148 201500 5160
rect 174044 5120 201500 5148
rect 174044 5108 174050 5120
rect 201494 5108 201500 5120
rect 201552 5108 201558 5160
rect 213914 5108 213920 5160
rect 213972 5148 213978 5160
rect 296070 5148 296076 5160
rect 213972 5120 296076 5148
rect 213972 5108 213978 5120
rect 296070 5108 296076 5120
rect 296128 5108 296134 5160
rect 306374 5108 306380 5160
rect 306432 5148 306438 5160
rect 523034 5148 523040 5160
rect 306432 5120 523040 5148
rect 306432 5108 306438 5120
rect 523034 5108 523040 5120
rect 523092 5108 523098 5160
rect 21818 5040 21824 5092
rect 21876 5080 21882 5092
rect 100846 5080 100852 5092
rect 21876 5052 100852 5080
rect 21876 5040 21882 5052
rect 100846 5040 100852 5052
rect 100904 5040 100910 5092
rect 118602 5040 118608 5092
rect 118660 5080 118666 5092
rect 139486 5080 139492 5092
rect 118660 5052 139492 5080
rect 118660 5040 118666 5052
rect 139486 5040 139492 5052
rect 139544 5040 139550 5092
rect 175366 5040 175372 5092
rect 175424 5080 175430 5092
rect 205082 5080 205088 5092
rect 175424 5052 205088 5080
rect 175424 5040 175430 5052
rect 205082 5040 205088 5052
rect 205140 5040 205146 5092
rect 211154 5040 211160 5092
rect 211212 5080 211218 5092
rect 292574 5080 292580 5092
rect 211212 5052 292580 5080
rect 211212 5040 211218 5052
rect 292574 5040 292580 5052
rect 292632 5040 292638 5092
rect 307754 5040 307760 5092
rect 307812 5080 307818 5092
rect 526622 5080 526628 5092
rect 307812 5052 526628 5080
rect 307812 5040 307818 5052
rect 526622 5040 526628 5052
rect 526680 5040 526686 5092
rect 17034 4972 17040 5024
rect 17092 5012 17098 5024
rect 98178 5012 98184 5024
rect 17092 4984 98184 5012
rect 17092 4972 17098 4984
rect 98178 4972 98184 4984
rect 98236 4972 98242 5024
rect 104526 4972 104532 5024
rect 104584 5012 104590 5024
rect 133966 5012 133972 5024
rect 104584 4984 133972 5012
rect 104584 4972 104590 4984
rect 133966 4972 133972 4984
rect 134024 4972 134030 5024
rect 176838 4972 176844 5024
rect 176896 5012 176902 5024
rect 208578 5012 208584 5024
rect 176896 4984 208584 5012
rect 176896 4972 176902 4984
rect 208578 4972 208584 4984
rect 208636 4972 208642 5024
rect 215294 4972 215300 5024
rect 215352 5012 215358 5024
rect 299658 5012 299664 5024
rect 215352 4984 299664 5012
rect 215352 4972 215358 4984
rect 299658 4972 299664 4984
rect 299716 4972 299722 5024
rect 309134 4972 309140 5024
rect 309192 5012 309198 5024
rect 530118 5012 530124 5024
rect 309192 4984 530124 5012
rect 309192 4972 309198 4984
rect 530118 4972 530124 4984
rect 530176 4972 530182 5024
rect 12342 4904 12348 4956
rect 12400 4944 12406 4956
rect 96614 4944 96620 4956
rect 12400 4916 96620 4944
rect 12400 4904 12406 4916
rect 96614 4904 96620 4916
rect 96672 4904 96678 4956
rect 101030 4904 101036 4956
rect 101088 4944 101094 4956
rect 132678 4944 132684 4956
rect 101088 4916 132684 4944
rect 101088 4904 101094 4916
rect 132678 4904 132684 4916
rect 132736 4904 132742 4956
rect 178218 4904 178224 4956
rect 178276 4944 178282 4956
rect 209774 4944 209780 4956
rect 178276 4916 209780 4944
rect 178276 4904 178282 4916
rect 209774 4904 209780 4916
rect 209832 4904 209838 4956
rect 216674 4904 216680 4956
rect 216732 4944 216738 4956
rect 303154 4944 303160 4956
rect 216732 4916 303160 4944
rect 216732 4904 216738 4916
rect 303154 4904 303160 4916
rect 303212 4904 303218 4956
rect 310514 4904 310520 4956
rect 310572 4944 310578 4956
rect 533706 4944 533712 4956
rect 310572 4916 533712 4944
rect 310572 4904 310578 4916
rect 533706 4904 533712 4916
rect 533764 4904 533770 4956
rect 8754 4836 8760 4888
rect 8812 4876 8818 4888
rect 95326 4876 95332 4888
rect 8812 4848 95332 4876
rect 8812 4836 8818 4848
rect 95326 4836 95332 4848
rect 95384 4836 95390 4888
rect 97442 4836 97448 4888
rect 97500 4876 97506 4888
rect 131206 4876 131212 4888
rect 97500 4848 131212 4876
rect 97500 4836 97506 4848
rect 131206 4836 131212 4848
rect 131264 4836 131270 4888
rect 178126 4836 178132 4888
rect 178184 4876 178190 4888
rect 212166 4876 212172 4888
rect 178184 4848 212172 4876
rect 178184 4836 178190 4848
rect 212166 4836 212172 4848
rect 212224 4836 212230 4888
rect 218146 4836 218152 4888
rect 218204 4876 218210 4888
rect 306742 4876 306748 4888
rect 218204 4848 306748 4876
rect 218204 4836 218210 4848
rect 306742 4836 306748 4848
rect 306800 4836 306806 4888
rect 314654 4836 314660 4888
rect 314712 4876 314718 4888
rect 540790 4876 540796 4888
rect 314712 4848 540796 4876
rect 314712 4836 314718 4848
rect 540790 4836 540796 4848
rect 540848 4836 540854 4888
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 92566 4808 92572 4820
rect 4120 4780 92572 4808
rect 4120 4768 4126 4780
rect 92566 4768 92572 4780
rect 92624 4768 92630 4820
rect 93946 4768 93952 4820
rect 94004 4808 94010 4820
rect 129826 4808 129832 4820
rect 94004 4780 129832 4808
rect 94004 4768 94010 4780
rect 129826 4768 129832 4780
rect 129884 4768 129890 4820
rect 180794 4768 180800 4820
rect 180852 4808 180858 4820
rect 216858 4808 216864 4820
rect 180852 4780 216864 4808
rect 180852 4768 180858 4780
rect 216858 4768 216864 4780
rect 216916 4768 216922 4820
rect 220814 4768 220820 4820
rect 220872 4808 220878 4820
rect 313826 4808 313832 4820
rect 220872 4780 313832 4808
rect 220872 4768 220878 4780
rect 313826 4768 313832 4780
rect 313884 4768 313890 4820
rect 316034 4768 316040 4820
rect 316092 4808 316098 4820
rect 544378 4808 544384 4820
rect 316092 4780 544384 4808
rect 316092 4768 316098 4780
rect 544378 4768 544384 4780
rect 544436 4768 544442 4820
rect 83274 4700 83280 4752
rect 83332 4740 83338 4752
rect 125686 4740 125692 4752
rect 83332 4712 125692 4740
rect 83332 4700 83338 4712
rect 125686 4700 125692 4712
rect 125744 4700 125750 4752
rect 193306 4700 193312 4752
rect 193364 4740 193370 4752
rect 246390 4740 246396 4752
rect 193364 4712 246396 4740
rect 193364 4700 193370 4712
rect 246390 4700 246396 4712
rect 246448 4700 246454 4752
rect 257430 4700 257436 4752
rect 257488 4740 257494 4752
rect 286594 4740 286600 4752
rect 257488 4712 286600 4740
rect 257488 4700 257494 4712
rect 286594 4700 286600 4712
rect 286652 4700 286658 4752
rect 298094 4700 298100 4752
rect 298152 4740 298158 4752
rect 501782 4740 501788 4752
rect 298152 4712 501788 4740
rect 298152 4700 298158 4712
rect 501782 4700 501788 4712
rect 501840 4700 501846 4752
rect 86862 4632 86868 4684
rect 86920 4672 86926 4684
rect 126974 4672 126980 4684
rect 86920 4644 126980 4672
rect 86920 4632 86926 4644
rect 126974 4632 126980 4644
rect 127032 4632 127038 4684
rect 191926 4632 191932 4684
rect 191984 4672 191990 4684
rect 242894 4672 242900 4684
rect 191984 4644 242900 4672
rect 191984 4632 191990 4644
rect 242894 4632 242900 4644
rect 242952 4632 242958 4684
rect 296714 4632 296720 4684
rect 296772 4672 296778 4684
rect 498194 4672 498200 4684
rect 296772 4644 498200 4672
rect 296772 4632 296778 4644
rect 498194 4632 498200 4644
rect 498252 4632 498258 4684
rect 90358 4564 90364 4616
rect 90416 4604 90422 4616
rect 128446 4604 128452 4616
rect 90416 4576 128452 4604
rect 90416 4564 90422 4576
rect 128446 4564 128452 4576
rect 128504 4564 128510 4616
rect 183646 4564 183652 4616
rect 183704 4604 183710 4616
rect 221734 4604 221740 4616
rect 183704 4576 221740 4604
rect 183704 4564 183710 4576
rect 221734 4564 221740 4576
rect 221792 4564 221798 4616
rect 243538 4564 243544 4616
rect 243596 4604 243602 4616
rect 320910 4604 320916 4616
rect 243596 4576 320916 4604
rect 243596 4564 243602 4576
rect 320910 4564 320916 4576
rect 320968 4564 320974 4616
rect 115198 4496 115204 4548
rect 115256 4536 115262 4548
rect 135346 4536 135352 4548
rect 115256 4508 135352 4536
rect 115256 4496 115262 4508
rect 135346 4496 135352 4508
rect 135404 4496 135410 4548
rect 182358 4496 182364 4548
rect 182416 4536 182422 4548
rect 219250 4536 219256 4548
rect 182416 4508 219256 4536
rect 182416 4496 182422 4508
rect 219250 4496 219256 4508
rect 219308 4496 219314 4548
rect 242158 4496 242164 4548
rect 242216 4536 242222 4548
rect 317322 4536 317328 4548
rect 242216 4508 317328 4536
rect 242216 4496 242222 4508
rect 317322 4496 317328 4508
rect 317380 4496 317386 4548
rect 190546 4428 190552 4480
rect 190604 4468 190610 4480
rect 222470 4468 222476 4480
rect 190604 4440 222476 4468
rect 190604 4428 190610 4440
rect 222470 4428 222476 4440
rect 222528 4428 222534 4480
rect 243446 4156 243452 4208
rect 243504 4196 243510 4208
rect 243504 4168 243768 4196
rect 243504 4156 243510 4168
rect 67910 4088 67916 4140
rect 67968 4128 67974 4140
rect 118694 4128 118700 4140
rect 67968 4100 118700 4128
rect 67968 4088 67974 4100
rect 118694 4088 118700 4100
rect 118752 4088 118758 4140
rect 130562 4088 130568 4140
rect 130620 4128 130626 4140
rect 144914 4128 144920 4140
rect 130620 4100 144920 4128
rect 130620 4088 130626 4100
rect 144914 4088 144920 4100
rect 144972 4088 144978 4140
rect 158990 4088 158996 4140
rect 159048 4128 159054 4140
rect 163682 4128 163688 4140
rect 159048 4100 163688 4128
rect 159048 4088 159054 4100
rect 163682 4088 163688 4100
rect 163740 4088 163746 4140
rect 172514 4088 172520 4140
rect 172572 4128 172578 4140
rect 195606 4128 195612 4140
rect 172572 4100 195612 4128
rect 172572 4088 172578 4100
rect 195606 4088 195612 4100
rect 195664 4088 195670 4140
rect 199378 4088 199384 4140
rect 199436 4128 199442 4140
rect 202690 4128 202696 4140
rect 199436 4100 202696 4128
rect 199436 4088 199442 4100
rect 202690 4088 202696 4100
rect 202748 4088 202754 4140
rect 220078 4088 220084 4140
rect 220136 4128 220142 4140
rect 220538 4128 220544 4140
rect 220136 4100 220544 4128
rect 220136 4088 220142 4100
rect 220538 4088 220544 4100
rect 220596 4088 220602 4140
rect 232498 4088 232504 4140
rect 232556 4128 232562 4140
rect 243630 4128 243636 4140
rect 232556 4100 243636 4128
rect 232556 4088 232562 4100
rect 243630 4088 243636 4100
rect 243688 4088 243694 4140
rect 243740 4128 243768 4168
rect 268838 4128 268844 4140
rect 243740 4100 268844 4128
rect 268838 4088 268844 4100
rect 268896 4088 268902 4140
rect 277394 4088 277400 4140
rect 277452 4128 277458 4140
rect 450906 4128 450912 4140
rect 277452 4100 450912 4128
rect 277452 4088 277458 4100
rect 450906 4088 450912 4100
rect 450964 4088 450970 4140
rect 60826 4020 60832 4072
rect 60884 4060 60890 4072
rect 116026 4060 116032 4072
rect 60884 4032 116032 4060
rect 60884 4020 60890 4032
rect 116026 4020 116032 4032
rect 116084 4020 116090 4072
rect 129366 4020 129372 4072
rect 129424 4060 129430 4072
rect 145006 4060 145012 4072
rect 129424 4032 145012 4060
rect 129424 4020 129430 4032
rect 145006 4020 145012 4032
rect 145064 4020 145070 4072
rect 160094 4020 160100 4072
rect 160152 4060 160158 4072
rect 168374 4060 168380 4072
rect 160152 4032 168380 4060
rect 160152 4020 160158 4032
rect 168374 4020 168380 4032
rect 168432 4020 168438 4072
rect 173894 4020 173900 4072
rect 173952 4060 173958 4072
rect 199102 4060 199108 4072
rect 173952 4032 199108 4060
rect 173952 4020 173958 4032
rect 199102 4020 199108 4032
rect 199160 4020 199166 4072
rect 215938 4020 215944 4072
rect 215996 4060 216002 4072
rect 225138 4060 225144 4072
rect 215996 4032 225144 4060
rect 215996 4020 216002 4032
rect 225138 4020 225144 4032
rect 225196 4020 225202 4072
rect 226978 4020 226984 4072
rect 227036 4060 227042 4072
rect 264146 4060 264152 4072
rect 227036 4032 264152 4060
rect 227036 4020 227042 4032
rect 264146 4020 264152 4032
rect 264204 4020 264210 4072
rect 278774 4020 278780 4072
rect 278832 4060 278838 4072
rect 454494 4060 454500 4072
rect 278832 4032 454500 4060
rect 278832 4020 278838 4032
rect 454494 4020 454500 4032
rect 454552 4020 454558 4072
rect 53742 3952 53748 4004
rect 53800 3992 53806 4004
rect 113174 3992 113180 4004
rect 53800 3964 113180 3992
rect 53800 3952 53806 3964
rect 113174 3952 113180 3964
rect 113232 3952 113238 4004
rect 126974 3952 126980 4004
rect 127032 3992 127038 4004
rect 143626 3992 143632 4004
rect 127032 3964 143632 3992
rect 127032 3952 127038 3964
rect 143626 3952 143632 3964
rect 143684 3952 143690 4004
rect 161566 3952 161572 4004
rect 161624 3992 161630 4004
rect 171962 3992 171968 4004
rect 161624 3964 171968 3992
rect 161624 3952 161630 3964
rect 171962 3952 171968 3964
rect 172020 3952 172026 4004
rect 176746 3952 176752 4004
rect 176804 3992 176810 4004
rect 206186 3992 206192 4004
rect 176804 3964 206192 3992
rect 176804 3952 176810 3964
rect 206186 3952 206192 3964
rect 206244 3952 206250 4004
rect 216766 3952 216772 4004
rect 216824 3992 216830 4004
rect 228726 3992 228732 4004
rect 216824 3964 228732 3992
rect 216824 3952 216830 3964
rect 228726 3952 228732 3964
rect 228784 3952 228790 4004
rect 229738 3952 229744 4004
rect 229796 3992 229802 4004
rect 267734 3992 267740 4004
rect 229796 3964 267740 3992
rect 229796 3952 229802 3964
rect 267734 3952 267740 3964
rect 267792 3952 267798 4004
rect 280154 3952 280160 4004
rect 280212 3992 280218 4004
rect 458082 3992 458088 4004
rect 280212 3964 458088 3992
rect 280212 3952 280218 3964
rect 458082 3952 458088 3964
rect 458140 3952 458146 4004
rect 46658 3884 46664 3936
rect 46716 3924 46722 3936
rect 110414 3924 110420 3936
rect 46716 3896 110420 3924
rect 46716 3884 46722 3896
rect 110414 3884 110420 3896
rect 110472 3884 110478 3936
rect 125870 3884 125876 3936
rect 125928 3924 125934 3936
rect 143718 3924 143724 3936
rect 125928 3896 143724 3924
rect 125928 3884 125934 3896
rect 143718 3884 143724 3896
rect 143776 3884 143782 3936
rect 162854 3884 162860 3936
rect 162912 3924 162918 3936
rect 173158 3924 173164 3936
rect 162912 3896 173164 3924
rect 162912 3884 162918 3896
rect 173158 3884 173164 3896
rect 173216 3884 173222 3936
rect 179414 3884 179420 3936
rect 179472 3924 179478 3936
rect 213362 3924 213368 3936
rect 179472 3896 213368 3924
rect 179472 3884 179478 3896
rect 213362 3884 213368 3896
rect 213420 3884 213426 3936
rect 218054 3884 218060 3936
rect 218112 3924 218118 3936
rect 232222 3924 232228 3936
rect 218112 3896 232228 3924
rect 218112 3884 218118 3896
rect 232222 3884 232228 3896
rect 232280 3884 232286 3936
rect 235258 3884 235264 3936
rect 235316 3924 235322 3936
rect 235316 3896 243584 3924
rect 235316 3884 235322 3896
rect 39574 3816 39580 3868
rect 39632 3856 39638 3868
rect 107654 3856 107660 3868
rect 39632 3828 107660 3856
rect 39632 3816 39638 3828
rect 107654 3816 107660 3828
rect 107712 3816 107718 3868
rect 123478 3816 123484 3868
rect 123536 3856 123542 3868
rect 142246 3856 142252 3868
rect 123536 3828 142252 3856
rect 123536 3816 123542 3828
rect 142246 3816 142252 3828
rect 142304 3816 142310 3868
rect 162946 3816 162952 3868
rect 163004 3856 163010 3868
rect 174262 3856 174268 3868
rect 163004 3828 174268 3856
rect 163004 3816 163010 3828
rect 174262 3816 174268 3828
rect 174320 3816 174326 3868
rect 182266 3816 182272 3868
rect 182324 3856 182330 3868
rect 220446 3856 220452 3868
rect 182324 3828 220452 3856
rect 182324 3816 182330 3828
rect 220446 3816 220452 3828
rect 220504 3816 220510 3868
rect 220538 3816 220544 3868
rect 220596 3856 220602 3868
rect 235810 3856 235816 3868
rect 220596 3828 235816 3856
rect 220596 3816 220602 3828
rect 235810 3816 235816 3828
rect 235868 3816 235874 3868
rect 237374 3816 237380 3868
rect 237432 3856 237438 3868
rect 243446 3856 243452 3868
rect 237432 3828 243452 3856
rect 237432 3816 237438 3828
rect 243446 3816 243452 3828
rect 243504 3816 243510 3868
rect 243556 3856 243584 3896
rect 243630 3884 243636 3936
rect 243688 3924 243694 3936
rect 274818 3924 274824 3936
rect 243688 3896 274824 3924
rect 243688 3884 243694 3896
rect 274818 3884 274824 3896
rect 274876 3884 274882 3936
rect 281534 3884 281540 3936
rect 281592 3924 281598 3936
rect 461578 3924 461584 3936
rect 281592 3896 461584 3924
rect 281592 3884 281598 3896
rect 461578 3884 461584 3896
rect 461636 3884 461642 3936
rect 278314 3856 278320 3868
rect 243556 3828 278320 3856
rect 278314 3816 278320 3828
rect 278372 3816 278378 3868
rect 282914 3816 282920 3868
rect 282972 3856 282978 3868
rect 465166 3856 465172 3868
rect 282972 3828 465172 3856
rect 282972 3816 282978 3828
rect 465166 3816 465172 3828
rect 465224 3816 465230 3868
rect 32398 3748 32404 3800
rect 32456 3788 32462 3800
rect 104986 3788 104992 3800
rect 32456 3760 104992 3788
rect 32456 3748 32462 3760
rect 104986 3748 104992 3760
rect 105044 3748 105050 3800
rect 121086 3748 121092 3800
rect 121144 3788 121150 3800
rect 140774 3788 140780 3800
rect 121144 3760 140780 3788
rect 121144 3748 121150 3760
rect 140774 3748 140780 3760
rect 140832 3748 140838 3800
rect 142430 3748 142436 3800
rect 142488 3788 142494 3800
rect 150618 3788 150624 3800
rect 142488 3760 150624 3788
rect 142488 3748 142494 3760
rect 150618 3748 150624 3760
rect 150676 3748 150682 3800
rect 164234 3748 164240 3800
rect 164292 3788 164298 3800
rect 176654 3788 176660 3800
rect 164292 3760 176660 3788
rect 164292 3748 164298 3760
rect 176654 3748 176660 3760
rect 176712 3748 176718 3800
rect 186314 3748 186320 3800
rect 186372 3788 186378 3800
rect 231026 3788 231032 3800
rect 186372 3760 231032 3788
rect 186372 3748 186378 3760
rect 231026 3748 231032 3760
rect 231084 3748 231090 3800
rect 233878 3748 233884 3800
rect 233936 3788 233942 3800
rect 281902 3788 281908 3800
rect 233936 3760 281908 3788
rect 233936 3748 233942 3760
rect 281902 3748 281908 3760
rect 281960 3748 281966 3800
rect 284478 3748 284484 3800
rect 284536 3788 284542 3800
rect 468662 3788 468668 3800
rect 284536 3760 468668 3788
rect 284536 3748 284542 3760
rect 468662 3748 468668 3760
rect 468720 3748 468726 3800
rect 24210 3680 24216 3732
rect 24268 3720 24274 3732
rect 100754 3720 100760 3732
rect 24268 3692 100760 3720
rect 24268 3680 24274 3692
rect 100754 3680 100760 3692
rect 100812 3680 100818 3732
rect 111610 3680 111616 3732
rect 111668 3720 111674 3732
rect 117222 3720 117228 3732
rect 111668 3692 117228 3720
rect 111668 3680 111674 3692
rect 117222 3680 117228 3692
rect 117280 3680 117286 3732
rect 119890 3680 119896 3732
rect 119948 3720 119954 3732
rect 140866 3720 140872 3732
rect 119948 3692 140872 3720
rect 119948 3680 119954 3692
rect 140866 3680 140872 3692
rect 140924 3680 140930 3732
rect 149146 3720 149152 3732
rect 142126 3692 149152 3720
rect 15930 3612 15936 3664
rect 15988 3652 15994 3664
rect 97994 3652 98000 3664
rect 15988 3624 98000 3652
rect 15988 3612 15994 3624
rect 97994 3612 98000 3624
rect 98052 3612 98058 3664
rect 118786 3612 118792 3664
rect 118844 3652 118850 3664
rect 140958 3652 140964 3664
rect 118844 3624 140964 3652
rect 118844 3612 118850 3624
rect 140958 3612 140964 3624
rect 141016 3612 141022 3664
rect 141234 3612 141240 3664
rect 141292 3652 141298 3664
rect 142126 3652 142154 3692
rect 149146 3680 149152 3692
rect 149204 3680 149210 3732
rect 157518 3680 157524 3732
rect 157576 3720 157582 3732
rect 161290 3720 161296 3732
rect 157576 3692 161296 3720
rect 157576 3680 157582 3692
rect 161290 3680 161296 3692
rect 161348 3680 161354 3732
rect 165706 3680 165712 3732
rect 165764 3720 165770 3732
rect 180242 3720 180248 3732
rect 165764 3692 180248 3720
rect 165764 3680 165770 3692
rect 180242 3680 180248 3692
rect 180300 3680 180306 3732
rect 189166 3680 189172 3732
rect 189224 3720 189230 3732
rect 238110 3720 238116 3732
rect 189224 3692 238116 3720
rect 189224 3680 189230 3692
rect 238110 3680 238116 3692
rect 238168 3680 238174 3732
rect 240134 3680 240140 3732
rect 240192 3720 240198 3732
rect 272426 3720 272432 3732
rect 240192 3692 272432 3720
rect 240192 3680 240198 3692
rect 272426 3680 272432 3692
rect 272484 3680 272490 3732
rect 285674 3680 285680 3732
rect 285732 3720 285738 3732
rect 472250 3720 472256 3732
rect 285732 3692 472256 3720
rect 285732 3680 285738 3692
rect 472250 3680 472256 3692
rect 472308 3680 472314 3732
rect 147858 3652 147864 3664
rect 141292 3624 142154 3652
rect 145024 3624 147864 3652
rect 141292 3612 141298 3624
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 95418 3584 95424 3596
rect 11204 3556 95424 3584
rect 11204 3544 11210 3556
rect 95418 3544 95424 3556
rect 95476 3544 95482 3596
rect 102226 3544 102232 3596
rect 102284 3584 102290 3596
rect 108298 3584 108304 3596
rect 102284 3556 108304 3584
rect 102284 3544 102290 3556
rect 108298 3544 108304 3556
rect 108356 3544 108362 3596
rect 114002 3544 114008 3596
rect 114060 3584 114066 3596
rect 138106 3584 138112 3596
rect 114060 3556 138112 3584
rect 114060 3544 114066 3556
rect 138106 3544 138112 3556
rect 138164 3544 138170 3596
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 98086 3516 98092 3528
rect 14792 3488 98092 3516
rect 14792 3476 14798 3488
rect 98086 3476 98092 3488
rect 98144 3476 98150 3528
rect 103330 3476 103336 3528
rect 103388 3516 103394 3528
rect 134058 3516 134064 3528
rect 103388 3488 134064 3516
rect 103388 3476 103394 3488
rect 134058 3476 134064 3488
rect 134116 3476 134122 3528
rect 135254 3476 135260 3528
rect 135312 3516 135318 3528
rect 145024 3516 145052 3624
rect 147858 3612 147864 3624
rect 147916 3612 147922 3664
rect 157426 3612 157432 3664
rect 157484 3652 157490 3664
rect 160094 3652 160100 3664
rect 157484 3624 160100 3652
rect 157484 3612 157490 3624
rect 160094 3612 160100 3624
rect 160152 3612 160158 3664
rect 165614 3612 165620 3664
rect 165672 3652 165678 3664
rect 181438 3652 181444 3664
rect 165672 3624 181444 3652
rect 165672 3612 165678 3624
rect 181438 3612 181444 3624
rect 181496 3612 181502 3664
rect 190454 3612 190460 3664
rect 190512 3652 190518 3664
rect 241698 3652 241704 3664
rect 190512 3624 241704 3652
rect 190512 3612 190518 3624
rect 241698 3612 241704 3624
rect 241756 3612 241762 3664
rect 249794 3612 249800 3664
rect 249852 3652 249858 3664
rect 279510 3652 279516 3664
rect 249852 3624 279516 3652
rect 249852 3612 249858 3624
rect 279510 3612 279516 3624
rect 279568 3612 279574 3664
rect 287054 3612 287060 3664
rect 287112 3652 287118 3664
rect 475746 3652 475752 3664
rect 287112 3624 475752 3652
rect 287112 3612 287118 3624
rect 475746 3612 475752 3624
rect 475804 3612 475810 3664
rect 146478 3544 146484 3596
rect 146536 3544 146542 3596
rect 158806 3544 158812 3596
rect 158864 3544 158870 3596
rect 166994 3544 167000 3596
rect 167052 3584 167058 3596
rect 184934 3584 184940 3596
rect 167052 3556 184940 3584
rect 167052 3544 167058 3556
rect 184934 3544 184940 3556
rect 184992 3544 184998 3596
rect 191834 3544 191840 3596
rect 191892 3584 191898 3596
rect 245194 3584 245200 3596
rect 191892 3556 245200 3584
rect 191892 3544 191898 3556
rect 245194 3544 245200 3556
rect 245252 3544 245258 3596
rect 247678 3544 247684 3596
rect 247736 3584 247742 3596
rect 276014 3584 276020 3596
rect 247736 3556 276020 3584
rect 247736 3544 247742 3556
rect 276014 3544 276020 3556
rect 276072 3544 276078 3596
rect 331214 3544 331220 3596
rect 331272 3584 331278 3596
rect 582190 3584 582196 3596
rect 331272 3556 582196 3584
rect 331272 3544 331278 3556
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 135312 3488 145052 3516
rect 135312 3476 135318 3488
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 93854 3448 93860 3460
rect 6512 3420 93860 3448
rect 6512 3408 6518 3420
rect 93854 3408 93860 3420
rect 93912 3408 93918 3460
rect 96246 3408 96252 3460
rect 96304 3448 96310 3460
rect 131114 3448 131120 3460
rect 96304 3420 131120 3448
rect 96304 3408 96310 3420
rect 131114 3408 131120 3420
rect 131172 3408 131178 3460
rect 132954 3408 132960 3460
rect 133012 3448 133018 3460
rect 146496 3448 146524 3544
rect 153010 3476 153016 3528
rect 153068 3516 153074 3528
rect 154666 3516 154672 3528
rect 153068 3488 154672 3516
rect 153068 3476 153074 3488
rect 154666 3476 154672 3488
rect 154724 3476 154730 3528
rect 155954 3476 155960 3528
rect 156012 3516 156018 3528
rect 156230 3516 156236 3528
rect 156012 3488 156236 3516
rect 156012 3476 156018 3488
rect 156230 3476 156236 3488
rect 156288 3476 156294 3528
rect 158824 3516 158852 3544
rect 164510 3516 164516 3528
rect 158824 3488 164516 3516
rect 164510 3476 164516 3488
rect 164568 3476 164574 3528
rect 164878 3476 164884 3528
rect 164936 3516 164942 3528
rect 166074 3516 166080 3528
rect 164936 3488 166080 3516
rect 164936 3476 164942 3488
rect 166074 3476 166080 3488
rect 166132 3476 166138 3528
rect 168466 3476 168472 3528
rect 168524 3516 168530 3528
rect 188522 3516 188528 3528
rect 168524 3488 188528 3516
rect 168524 3476 168530 3488
rect 188522 3476 188528 3488
rect 188580 3476 188586 3528
rect 194594 3476 194600 3528
rect 194652 3516 194658 3528
rect 252370 3516 252376 3528
rect 194652 3488 252376 3516
rect 194652 3476 194658 3488
rect 252370 3476 252376 3488
rect 252428 3476 252434 3528
rect 258074 3476 258080 3528
rect 258132 3516 258138 3528
rect 266538 3516 266544 3528
rect 258132 3488 266544 3516
rect 258132 3476 258138 3488
rect 266538 3476 266544 3488
rect 266596 3476 266602 3528
rect 288434 3476 288440 3528
rect 288492 3516 288498 3528
rect 479334 3516 479340 3528
rect 288492 3488 479340 3516
rect 288492 3476 288498 3488
rect 479334 3476 479340 3488
rect 479392 3476 479398 3528
rect 489914 3476 489920 3528
rect 489972 3516 489978 3528
rect 490742 3516 490748 3528
rect 489972 3488 490748 3516
rect 489972 3476 489978 3488
rect 490742 3476 490748 3488
rect 490800 3476 490806 3528
rect 531314 3476 531320 3528
rect 531372 3516 531378 3528
rect 532142 3516 532148 3528
rect 531372 3488 532148 3516
rect 531372 3476 531378 3488
rect 532142 3476 532148 3488
rect 532200 3476 532206 3528
rect 556154 3476 556160 3528
rect 556212 3516 556218 3528
rect 556982 3516 556988 3528
rect 556212 3488 556988 3516
rect 556212 3476 556218 3488
rect 556982 3476 556988 3488
rect 557040 3476 557046 3528
rect 133012 3420 146524 3448
rect 133012 3408 133018 3420
rect 160186 3408 160192 3460
rect 160244 3448 160250 3460
rect 167178 3448 167184 3460
rect 160244 3420 167184 3448
rect 160244 3408 160250 3420
rect 167178 3408 167184 3420
rect 167236 3408 167242 3460
rect 169846 3408 169852 3460
rect 169904 3448 169910 3460
rect 192018 3448 192024 3460
rect 169904 3420 192024 3448
rect 169904 3408 169910 3420
rect 192018 3408 192024 3420
rect 192076 3408 192082 3460
rect 198734 3408 198740 3460
rect 198792 3448 198798 3460
rect 259454 3448 259460 3460
rect 198792 3420 259460 3448
rect 198792 3408 198798 3420
rect 259454 3408 259460 3420
rect 259512 3408 259518 3460
rect 324406 3408 324412 3460
rect 324464 3448 324470 3460
rect 325602 3448 325608 3460
rect 324464 3420 325608 3448
rect 324464 3408 324470 3420
rect 325602 3408 325608 3420
rect 325660 3408 325666 3460
rect 332686 3408 332692 3460
rect 332744 3448 332750 3460
rect 333882 3448 333888 3460
rect 332744 3420 333888 3448
rect 332744 3408 332750 3420
rect 333882 3408 333888 3420
rect 333940 3408 333946 3460
rect 333974 3408 333980 3460
rect 334032 3448 334038 3460
rect 580994 3448 581000 3460
rect 334032 3420 581000 3448
rect 334032 3408 334038 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 19334 3340 19340 3392
rect 19392 3380 19398 3392
rect 20254 3380 20260 3392
rect 19392 3352 20260 3380
rect 19392 3340 19398 3352
rect 20254 3340 20260 3352
rect 20312 3340 20318 3392
rect 74994 3340 75000 3392
rect 75052 3380 75058 3392
rect 122834 3380 122840 3392
rect 75052 3352 122840 3380
rect 75052 3340 75058 3352
rect 122834 3340 122840 3352
rect 122892 3340 122898 3392
rect 131758 3340 131764 3392
rect 131816 3380 131822 3392
rect 145098 3380 145104 3392
rect 131816 3352 145104 3380
rect 131816 3340 131822 3352
rect 145098 3340 145104 3352
rect 145156 3340 145162 3392
rect 161658 3340 161664 3392
rect 161716 3380 161722 3392
rect 169570 3380 169576 3392
rect 161716 3352 169576 3380
rect 161716 3340 161722 3352
rect 169570 3340 169576 3352
rect 169628 3340 169634 3392
rect 206278 3340 206284 3392
rect 206336 3380 206342 3392
rect 207382 3380 207388 3392
rect 206336 3352 207388 3380
rect 206336 3340 206342 3352
rect 207382 3340 207388 3352
rect 207440 3340 207446 3392
rect 210418 3340 210424 3392
rect 210476 3380 210482 3392
rect 214466 3380 214472 3392
rect 210476 3352 214472 3380
rect 210476 3340 210482 3352
rect 214466 3340 214472 3352
rect 214524 3340 214530 3392
rect 225598 3340 225604 3392
rect 225656 3380 225662 3392
rect 253474 3380 253480 3392
rect 225656 3352 253480 3380
rect 225656 3340 225662 3352
rect 253474 3340 253480 3352
rect 253532 3340 253538 3392
rect 276106 3340 276112 3392
rect 276164 3380 276170 3392
rect 447410 3380 447416 3392
rect 276164 3352 447416 3380
rect 276164 3340 276170 3352
rect 447410 3340 447416 3352
rect 447468 3340 447474 3392
rect 448514 3340 448520 3392
rect 448572 3380 448578 3392
rect 449802 3380 449808 3392
rect 448572 3352 449808 3380
rect 448572 3340 448578 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 82078 3272 82084 3324
rect 82136 3312 82142 3324
rect 125594 3312 125600 3324
rect 82136 3284 125600 3312
rect 82136 3272 82142 3284
rect 125594 3272 125600 3284
rect 125652 3272 125658 3324
rect 136450 3272 136456 3324
rect 136508 3312 136514 3324
rect 147766 3312 147772 3324
rect 136508 3284 147772 3312
rect 136508 3272 136514 3284
rect 147766 3272 147772 3284
rect 147824 3272 147830 3324
rect 224218 3272 224224 3324
rect 224276 3312 224282 3324
rect 249978 3312 249984 3324
rect 224276 3284 249984 3312
rect 224276 3272 224282 3284
rect 249978 3272 249984 3284
rect 250036 3272 250042 3324
rect 274634 3272 274640 3324
rect 274692 3312 274698 3324
rect 443822 3312 443828 3324
rect 274692 3284 443828 3312
rect 274692 3272 274698 3284
rect 443822 3272 443828 3284
rect 443880 3272 443886 3324
rect 89162 3204 89168 3256
rect 89220 3244 89226 3256
rect 128354 3244 128360 3256
rect 89220 3216 128360 3244
rect 89220 3204 89226 3216
rect 128354 3204 128360 3216
rect 128412 3204 128418 3256
rect 134150 3204 134156 3256
rect 134208 3244 134214 3256
rect 146386 3244 146392 3256
rect 134208 3216 146392 3244
rect 134208 3204 134214 3216
rect 146386 3204 146392 3216
rect 146444 3204 146450 3256
rect 222470 3204 222476 3256
rect 222528 3244 222534 3256
rect 239306 3244 239312 3256
rect 222528 3216 239312 3244
rect 222528 3204 222534 3216
rect 239306 3204 239312 3216
rect 239364 3204 239370 3256
rect 273254 3204 273260 3256
rect 273312 3244 273318 3256
rect 440326 3244 440332 3256
rect 273312 3216 440332 3244
rect 273312 3204 273318 3216
rect 440326 3204 440332 3216
rect 440384 3204 440390 3256
rect 209038 3136 209044 3188
rect 209096 3176 209102 3188
rect 210970 3176 210976 3188
rect 209096 3148 210976 3176
rect 209096 3136 209102 3148
rect 210970 3136 210976 3148
rect 211028 3136 211034 3188
rect 211798 3136 211804 3188
rect 211856 3176 211862 3188
rect 218054 3176 218060 3188
rect 211856 3148 218060 3176
rect 211856 3136 211862 3148
rect 218054 3136 218060 3148
rect 218112 3136 218118 3188
rect 329834 3136 329840 3188
rect 329892 3176 329898 3188
rect 333974 3176 333980 3188
rect 329892 3148 333980 3176
rect 329892 3136 329898 3148
rect 333974 3136 333980 3148
rect 334032 3136 334038 3188
rect 349154 3136 349160 3188
rect 349212 3176 349218 3188
rect 350442 3176 350448 3188
rect 349212 3148 350448 3176
rect 349212 3136 349218 3148
rect 350442 3136 350448 3148
rect 350500 3136 350506 3188
rect 357434 3136 357440 3188
rect 357492 3176 357498 3188
rect 358722 3176 358728 3188
rect 357492 3148 358728 3176
rect 357492 3136 357498 3148
rect 358722 3136 358728 3148
rect 358780 3136 358786 3188
rect 365806 3136 365812 3188
rect 365864 3176 365870 3188
rect 367002 3176 367008 3188
rect 365864 3148 367008 3176
rect 365864 3136 365870 3148
rect 367002 3136 367008 3148
rect 367060 3136 367066 3188
rect 373994 3136 374000 3188
rect 374052 3176 374058 3188
rect 375282 3176 375288 3188
rect 374052 3148 375288 3176
rect 374052 3136 374058 3148
rect 375282 3136 375288 3148
rect 375340 3136 375346 3188
rect 382274 3136 382280 3188
rect 382332 3176 382338 3188
rect 383562 3176 383568 3188
rect 382332 3148 383568 3176
rect 382332 3136 382338 3148
rect 383562 3136 383568 3148
rect 383620 3136 383626 3188
rect 398834 3136 398840 3188
rect 398892 3176 398898 3188
rect 400122 3176 400128 3188
rect 398892 3148 400128 3176
rect 398892 3136 398898 3148
rect 400122 3136 400128 3148
rect 400180 3136 400186 3188
rect 407114 3136 407120 3188
rect 407172 3176 407178 3188
rect 408402 3176 408408 3188
rect 407172 3148 408408 3176
rect 407172 3136 407178 3148
rect 408402 3136 408408 3148
rect 408460 3136 408466 3188
rect 423766 3136 423772 3188
rect 423824 3176 423830 3188
rect 424962 3176 424968 3188
rect 423824 3148 424968 3176
rect 423824 3136 423830 3148
rect 424962 3136 424968 3148
rect 425020 3136 425026 3188
rect 431954 3136 431960 3188
rect 432012 3176 432018 3188
rect 433242 3176 433248 3188
rect 432012 3148 433248 3176
rect 432012 3136 432018 3148
rect 433242 3136 433248 3148
rect 433300 3136 433306 3188
rect 145926 3068 145932 3120
rect 145984 3108 145990 3120
rect 151906 3108 151912 3120
rect 145984 3080 151912 3108
rect 145984 3068 145990 3080
rect 151906 3068 151912 3080
rect 151964 3068 151970 3120
rect 128170 3000 128176 3052
rect 128228 3040 128234 3052
rect 128998 3040 129004 3052
rect 128228 3012 129004 3040
rect 128228 3000 128234 3012
rect 128998 3000 129004 3012
rect 129056 3000 129062 3052
rect 144730 3000 144736 3052
rect 144788 3040 144794 3052
rect 150526 3040 150532 3052
rect 144788 3012 150532 3040
rect 144788 3000 144794 3012
rect 150526 3000 150532 3012
rect 150584 3000 150590 3052
rect 213178 3000 213184 3052
rect 213236 3040 213242 3052
rect 221550 3040 221556 3052
rect 213236 3012 221556 3040
rect 213236 3000 213242 3012
rect 221550 3000 221556 3012
rect 221608 3000 221614 3052
rect 149514 2932 149520 2984
rect 149572 2972 149578 2984
rect 153378 2972 153384 2984
rect 149572 2944 153384 2972
rect 149572 2932 149578 2944
rect 153378 2932 153384 2944
rect 153436 2932 153442 2984
rect 108114 2796 108120 2848
rect 108172 2836 108178 2848
rect 115198 2836 115204 2848
rect 108172 2808 115204 2836
rect 108172 2796 108178 2808
rect 115198 2796 115204 2808
rect 115256 2796 115262 2848
rect 115290 2796 115296 2848
rect 115348 2836 115354 2848
rect 118602 2836 118608 2848
rect 115348 2808 118608 2836
rect 115348 2796 115354 2808
rect 118602 2796 118608 2808
rect 118660 2796 118666 2848
rect 221734 2796 221740 2848
rect 221792 2836 221798 2848
rect 223942 2836 223948 2848
rect 221792 2808 223948 2836
rect 221792 2796 221798 2808
rect 223942 2796 223948 2808
rect 224000 2796 224006 2848
<< via1 >>
rect 137836 700952 137888 701004
rect 227720 700952 227772 701004
rect 208400 700884 208452 700936
rect 332508 700884 332560 700936
rect 209780 700816 209832 700868
rect 348792 700816 348844 700868
rect 89168 700748 89220 700800
rect 236000 700748 236052 700800
rect 72976 700680 73028 700732
rect 233240 700680 233292 700732
rect 201500 700612 201552 700664
rect 397460 700612 397512 700664
rect 204260 700544 204312 700596
rect 413652 700544 413704 700596
rect 24308 700476 24360 700528
rect 241520 700476 241572 700528
rect 8116 700408 8168 700460
rect 240140 700408 240192 700460
rect 197360 700340 197412 700392
rect 478512 700340 478564 700392
rect 191840 700272 191892 700324
rect 543464 700272 543516 700324
rect 154120 700204 154172 700256
rect 229100 700204 229152 700256
rect 202788 700136 202840 700188
rect 215944 700136 215996 700188
rect 216680 700136 216732 700188
rect 283840 700136 283892 700188
rect 218980 700068 219032 700120
rect 222200 700068 222252 700120
rect 183560 696940 183612 696992
rect 580172 696940 580224 696992
rect 266360 693472 266412 693524
rect 267648 693472 267700 693524
rect 3424 683204 3476 683256
rect 244280 683204 244332 683256
rect 184940 683136 184992 683188
rect 580172 683136 580224 683188
rect 3424 670760 3476 670812
rect 248420 670760 248472 670812
rect 180800 670692 180852 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 245660 656888 245712 656940
rect 176660 643084 176712 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 249800 632068 249852 632120
rect 178040 630640 178092 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 253940 618264 253992 618316
rect 173900 616836 173952 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 252560 605820 252612 605872
rect 169852 590656 169904 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 256700 579640 256752 579692
rect 172520 576852 172572 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 260840 565836 260892 565888
rect 168380 563048 168432 563100
rect 579804 563048 579856 563100
rect 3424 553392 3476 553444
rect 258080 553392 258132 553444
rect 164240 536800 164292 536852
rect 580172 536800 580224 536852
rect 3424 527144 3476 527196
rect 262220 527144 262272 527196
rect 165620 524424 165672 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 267740 514768 267792 514820
rect 161480 510620 161532 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 264980 500964 265032 501016
rect 157340 484372 157392 484424
rect 580172 484372 580224 484424
rect 3424 474716 3476 474768
rect 269120 474716 269172 474768
rect 160100 470568 160152 470620
rect 579988 470568 580040 470620
rect 3240 462340 3292 462392
rect 273260 462340 273312 462392
rect 155960 456764 156012 456816
rect 580172 456764 580224 456816
rect 3148 448536 3200 448588
rect 271880 448536 271932 448588
rect 151820 430584 151872 430636
rect 580172 430584 580224 430636
rect 3424 422288 3476 422340
rect 276020 422288 276072 422340
rect 153200 418140 153252 418192
rect 580172 418140 580224 418192
rect 3148 409844 3200 409896
rect 280160 409844 280212 409896
rect 149060 404336 149112 404388
rect 580172 404336 580224 404388
rect 3424 397468 3476 397520
rect 277400 397468 277452 397520
rect 144920 378156 144972 378208
rect 580172 378156 580224 378208
rect 3424 371220 3476 371272
rect 281540 371220 281592 371272
rect 147680 364352 147732 364404
rect 580172 364352 580224 364404
rect 3148 357416 3200 357468
rect 284944 357416 284996 357468
rect 143540 351908 143592 351960
rect 580172 351908 580224 351960
rect 109408 347760 109460 347812
rect 577688 347760 577740 347812
rect 215116 346332 215168 346384
rect 266360 346332 266412 346384
rect 169760 346264 169812 346316
rect 225604 346264 225656 346316
rect 213000 346196 213052 346248
rect 299480 346196 299532 346248
rect 104900 346128 104952 346180
rect 231952 346128 232004 346180
rect 206652 346060 206704 346112
rect 364340 346060 364392 346112
rect 40040 345992 40092 346044
rect 238300 345992 238352 346044
rect 200396 345924 200448 345976
rect 429200 345924 429252 345976
rect 196164 345856 196216 345908
rect 462320 345856 462372 345908
rect 194048 345788 194100 345840
rect 494060 345788 494112 345840
rect 189816 345720 189868 345772
rect 527180 345720 527232 345772
rect 187700 345652 187752 345704
rect 558920 345652 558972 345704
rect 219348 345584 219400 345636
rect 234620 345584 234672 345636
rect 3332 345040 3384 345092
rect 220820 345040 220872 345092
rect 215944 344496 215996 344548
rect 221464 344496 221516 344548
rect 220820 344428 220872 344480
rect 284576 344428 284628 344480
rect 284944 344428 284996 344480
rect 286692 344428 286744 344480
rect 126704 344360 126756 344412
rect 331956 344360 332008 344412
rect 114008 344292 114060 344344
rect 331864 344292 331916 344344
rect 90640 344224 90692 344276
rect 320364 344224 320416 344276
rect 3516 344156 3568 344208
rect 303528 344156 303580 344208
rect 3608 344088 3660 344140
rect 305644 344088 305696 344140
rect 4896 344020 4948 344072
rect 307760 344020 307812 344072
rect 3424 343952 3476 344004
rect 311992 343952 312044 344004
rect 4804 343884 4856 343936
rect 314108 343884 314160 343936
rect 92020 343816 92072 343868
rect 103520 343816 103572 343868
rect 105636 343816 105688 343868
rect 580264 343816 580316 343868
rect 92112 343748 92164 343800
rect 97172 343748 97224 343800
rect 101404 343748 101456 343800
rect 577596 343748 577648 343800
rect 95056 343680 95108 343732
rect 577504 343680 577556 343732
rect 93032 343612 93084 343664
rect 579620 343612 579672 343664
rect 90824 342728 90876 342780
rect 318248 342728 318300 342780
rect 90456 342660 90508 342712
rect 324596 342660 324648 342712
rect 3976 342592 4028 342644
rect 295156 342592 295208 342644
rect 3700 342524 3752 342576
rect 301412 342524 301464 342576
rect 124588 342456 124640 342508
rect 580816 342456 580868 342508
rect 122472 342388 122524 342440
rect 580632 342388 580684 342440
rect 118240 342320 118292 342372
rect 580540 342320 580592 342372
rect 111892 342252 111944 342304
rect 580448 342252 580500 342304
rect 135260 341776 135312 341828
rect 164792 341776 164844 341828
rect 90732 341436 90784 341488
rect 135260 341572 135312 341624
rect 135536 341572 135588 341624
rect 139952 341572 140004 341624
rect 3240 341368 3292 341420
rect 4068 341300 4120 341352
rect 135444 341504 135496 341556
rect 3332 341232 3384 341284
rect 135214 341436 135266 341488
rect 131120 341368 131172 341420
rect 135444 341368 135496 341420
rect 135536 341368 135588 341420
rect 3792 341164 3844 341216
rect 3884 341096 3936 341148
rect 137560 341368 137612 341420
rect 139584 341368 139636 341420
rect 139952 341368 140004 341420
rect 164148 341368 164200 341420
rect 164792 341368 164844 341420
rect 316040 341436 316092 341488
rect 288532 341368 288584 341420
rect 290556 341368 290608 341420
rect 292764 341368 292816 341420
rect 296904 341368 296956 341420
rect 299020 341368 299072 341420
rect 580080 341028 580132 341080
rect 580908 340960 580960 341012
rect 580172 340892 580224 340944
rect 331956 272552 332008 272604
rect 580080 272552 580132 272604
rect 331864 272484 331916 272536
rect 580908 272484 580960 272536
rect 2780 163752 2832 163804
rect 4896 163752 4948 163804
rect 2780 110712 2832 110764
rect 4804 110712 4856 110764
rect 161572 101804 161624 101856
rect 162768 101804 162820 101856
rect 241704 101736 241756 101788
rect 242624 101736 242676 101788
rect 329840 100920 329892 100972
rect 330760 100920 330812 100972
rect 325700 100784 325752 100836
rect 326344 100784 326396 100836
rect 70400 100648 70452 100700
rect 121368 100648 121420 100700
rect 171508 100648 171560 100700
rect 193220 100648 193272 100700
rect 194876 100648 194928 100700
rect 224224 100648 224276 100700
rect 577688 100648 577740 100700
rect 579988 100648 580040 100700
rect 63500 100580 63552 100632
rect 118424 100580 118476 100632
rect 129280 100580 129332 100632
rect 144736 100580 144788 100632
rect 146300 100580 146352 100632
rect 152556 100580 152608 100632
rect 177396 100580 177448 100632
rect 206284 100580 206336 100632
rect 208400 100580 208452 100632
rect 238024 100580 238076 100632
rect 56600 100512 56652 100564
rect 115572 100512 115624 100564
rect 125324 100512 125376 100564
rect 143264 100512 143316 100564
rect 157432 100512 157484 100564
rect 158720 100512 158772 100564
rect 172980 100512 173032 100564
rect 195980 100512 196032 100564
rect 196348 100512 196400 100564
rect 225512 100512 225564 100564
rect 49700 100444 49752 100496
rect 112628 100444 112680 100496
rect 117320 100444 117372 100496
rect 140320 100444 140372 100496
rect 156880 100444 156932 100496
rect 157340 100444 157392 100496
rect 174452 100444 174504 100496
rect 200120 100444 200172 100496
rect 206560 100444 206612 100496
rect 235356 100444 235408 100496
rect 264520 100444 264572 100496
rect 333244 100444 333296 100496
rect 42800 100376 42852 100428
rect 109684 100376 109736 100428
rect 121460 100376 121512 100428
rect 142344 100376 142396 100428
rect 170036 100376 170088 100428
rect 188988 100376 189040 100428
rect 189080 100376 189132 100428
rect 220084 100376 220136 100428
rect 224132 100376 224184 100428
rect 243360 100376 243412 100428
rect 288440 100376 288492 100428
rect 289360 100376 289412 100428
rect 331680 100376 331732 100428
rect 406384 100376 406436 100428
rect 35900 100308 35952 100360
rect 106740 100308 106792 100360
rect 115940 100308 115992 100360
rect 139860 100308 139912 100360
rect 158904 100308 158956 100360
rect 161480 100308 161532 100360
rect 167092 100308 167144 100360
rect 182180 100308 182232 100360
rect 183192 100308 183244 100360
rect 213184 100308 213236 100360
rect 222660 100308 222712 100360
rect 242164 100308 242216 100360
rect 252836 100308 252888 100360
rect 390560 100308 390612 100360
rect 27620 100240 27672 100292
rect 103888 100240 103940 100292
rect 108304 100240 108356 100292
rect 134064 100240 134116 100292
rect 137008 100240 137060 100292
rect 148600 100240 148652 100292
rect 151820 100240 151872 100292
rect 154488 100240 154540 100292
rect 181720 100240 181772 100292
rect 211804 100240 211856 100292
rect 212908 100240 212960 100292
rect 243636 100240 243688 100292
rect 255780 100240 255832 100292
rect 397460 100240 397512 100292
rect 19432 100172 19484 100224
rect 99932 100172 99984 100224
rect 111800 100172 111852 100224
rect 138388 100172 138440 100224
rect 148232 100172 148284 100224
rect 153016 100172 153068 100224
rect 167644 100172 167696 100224
rect 183560 100172 183612 100224
rect 184664 100172 184716 100224
rect 215944 100172 215996 100224
rect 224592 100172 224644 100224
rect 246304 100172 246356 100224
rect 258632 100172 258684 100224
rect 404360 100172 404412 100224
rect 24860 100104 24912 100156
rect 102416 100104 102468 100156
rect 106556 100104 106608 100156
rect 135996 100104 136048 100156
rect 139400 100104 139452 100156
rect 149612 100104 149664 100156
rect 164240 100104 164292 100156
rect 175280 100104 175332 100156
rect 175924 100104 175976 100156
rect 202880 100104 202932 100156
rect 205640 100104 205692 100156
rect 247684 100104 247736 100156
rect 261576 100104 261628 100156
rect 411260 100104 411312 100156
rect 19340 100036 19392 100088
rect 100392 100036 100444 100088
rect 110420 100036 110472 100088
rect 137468 100036 137520 100088
rect 165160 100036 165212 100088
rect 176936 100036 176988 100088
rect 180248 100036 180300 100088
rect 210424 100036 210476 100088
rect 211436 100036 211488 100088
rect 257344 100036 257396 100088
rect 267464 100036 267516 100088
rect 425060 100036 425112 100088
rect 9680 99968 9732 100020
rect 96068 99968 96120 100020
rect 104900 99968 104952 100020
rect 135444 99968 135496 100020
rect 138020 99968 138072 100020
rect 149152 99968 149204 100020
rect 150716 99968 150768 100020
rect 154028 99968 154080 100020
rect 160284 99968 160336 100020
rect 164884 99968 164936 100020
rect 165712 99968 165764 100020
rect 178040 99968 178092 100020
rect 178776 99968 178828 100020
rect 209044 99968 209096 100020
rect 209964 99968 210016 100020
rect 257436 99968 257488 100020
rect 270316 99968 270368 100020
rect 431960 99968 432012 100020
rect 77300 99900 77352 99952
rect 124312 99900 124364 99952
rect 165620 99900 165672 99952
rect 166632 99900 166684 99952
rect 175372 99900 175424 99952
rect 199384 99900 199436 99952
rect 205088 99900 205140 99952
rect 232504 99900 232556 99952
rect 305000 99900 305052 99952
rect 305920 99900 305972 99952
rect 92480 99832 92532 99884
rect 130108 99832 130160 99884
rect 168564 99832 168616 99884
rect 185308 99832 185360 99884
rect 202236 99832 202288 99884
rect 229744 99832 229796 99884
rect 99380 99764 99432 99816
rect 133052 99764 133104 99816
rect 208032 99764 208084 99816
rect 233884 99764 233936 99816
rect 93860 99696 93912 99748
rect 94596 99696 94648 99748
rect 200764 99696 200816 99748
rect 226892 99696 226944 99748
rect 285772 99628 285824 99680
rect 286876 99628 286928 99680
rect 143540 99560 143592 99612
rect 151084 99560 151136 99612
rect 162308 99492 162360 99544
rect 169760 99492 169812 99544
rect 248328 99424 248380 99476
rect 248972 99424 249024 99476
rect 168380 99220 168432 99272
rect 169576 99220 169628 99272
rect 287060 98608 287112 98660
rect 287888 98608 287940 98660
rect 158812 98472 158864 98524
rect 159824 98472 159876 98524
rect 249800 98200 249852 98252
rect 250352 98200 250404 98252
rect 133972 98132 134024 98184
rect 134984 98132 135036 98184
rect 185032 98064 185084 98116
rect 185676 98064 185728 98116
rect 229100 98064 229152 98116
rect 229928 98064 229980 98116
rect 110604 97996 110656 98048
rect 111616 97996 111668 98048
rect 127072 97996 127124 98048
rect 128176 97996 128228 98048
rect 131120 97996 131172 98048
rect 131580 97996 131632 98048
rect 186412 97996 186464 98048
rect 187608 97996 187660 98048
rect 203064 97996 203116 98048
rect 204168 97996 204220 98048
rect 225144 97996 225196 98048
rect 226064 97996 226116 98048
rect 226432 97996 226484 98048
rect 227536 97996 227588 98048
rect 251272 97996 251324 98048
rect 252376 97996 252428 98048
rect 254032 97996 254084 98048
rect 255228 97996 255280 98048
rect 284392 97996 284444 98048
rect 285404 97996 285456 98048
rect 292672 97996 292724 98048
rect 293684 97996 293736 98048
rect 294052 97996 294104 98048
rect 295156 97996 295208 98048
rect 295432 97996 295484 98048
rect 296628 97996 296680 98048
rect 317512 97996 317564 98048
rect 318524 97996 318576 98048
rect 318892 97996 318944 98048
rect 319996 97996 320048 98048
rect 320272 97996 320324 98048
rect 321468 97996 321520 98048
rect 3424 97928 3476 97980
rect 90824 97928 90876 97980
rect 91100 97928 91152 97980
rect 92204 97928 92256 97980
rect 92572 97928 92624 97980
rect 93584 97928 93636 97980
rect 100760 97928 100812 97980
rect 101864 97928 101916 97980
rect 102232 97928 102284 97980
rect 103336 97928 103388 97980
rect 103612 97928 103664 97980
rect 104808 97928 104860 97980
rect 107660 97928 107712 97980
rect 108212 97928 108264 97980
rect 110512 97928 110564 97980
rect 111156 97928 111208 97980
rect 113180 97928 113232 97980
rect 114100 97928 114152 97980
rect 118700 97928 118752 97980
rect 119896 97928 119948 97980
rect 120172 97928 120224 97980
rect 120908 97928 120960 97980
rect 126980 97928 127032 97980
rect 127716 97928 127768 97980
rect 131212 97928 131264 97980
rect 132040 97928 132092 97980
rect 140780 97928 140832 97980
rect 141792 97928 141844 97980
rect 143632 97928 143684 97980
rect 144276 97928 144328 97980
rect 144920 97928 144972 97980
rect 145748 97928 145800 97980
rect 146392 97928 146444 97980
rect 147220 97928 147272 97980
rect 160100 97928 160152 97980
rect 161296 97928 161348 97980
rect 169852 97928 169904 97980
rect 171048 97928 171100 97980
rect 178132 97928 178184 97980
rect 179328 97928 179380 97980
rect 185216 97928 185268 97980
rect 186136 97928 186188 97980
rect 186320 97928 186372 97980
rect 187056 97928 187108 97980
rect 189172 97928 189224 97980
rect 190000 97928 190052 97980
rect 190460 97928 190512 97980
rect 191472 97928 191524 97980
rect 191840 97928 191892 97980
rect 192944 97928 192996 97980
rect 194600 97928 194652 97980
rect 195888 97928 195940 97980
rect 202972 97928 203024 97980
rect 203616 97928 203668 97980
rect 208400 97928 208452 97980
rect 209504 97928 209556 97980
rect 209780 97928 209832 97980
rect 210976 97928 211028 97980
rect 211160 97928 211212 97980
rect 212448 97928 212500 97980
rect 224960 97928 225012 97980
rect 225604 97928 225656 97980
rect 226340 97928 226392 97980
rect 226984 97928 227036 97980
rect 227720 97928 227772 97980
rect 228456 97928 228508 97980
rect 230480 97928 230532 97980
rect 231400 97928 231452 97980
rect 233240 97928 233292 97980
rect 234344 97928 234396 97980
rect 234620 97928 234672 97980
rect 235816 97928 235868 97980
rect 241520 97928 241572 97980
rect 242072 97928 242124 97980
rect 242900 97928 242952 97980
rect 243544 97928 243596 97980
rect 244280 97928 244332 97980
rect 245016 97928 245068 97980
rect 248512 97928 248564 97980
rect 249432 97928 249484 97980
rect 251180 97928 251232 97980
rect 251824 97928 251876 97980
rect 253940 97928 253992 97980
rect 254768 97928 254820 97980
rect 258080 97928 258132 97980
rect 259184 97928 259236 97980
rect 259460 97928 259512 97980
rect 260656 97928 260708 97980
rect 260840 97928 260892 97980
rect 262036 97928 262088 97980
rect 262220 97928 262272 97980
rect 263508 97928 263560 97980
rect 266360 97928 266412 97980
rect 266912 97928 266964 97980
rect 267740 97928 267792 97980
rect 268384 97928 268436 97980
rect 269120 97928 269172 97980
rect 269856 97928 269908 97980
rect 270500 97928 270552 97980
rect 271328 97928 271380 97980
rect 271880 97928 271932 97980
rect 272800 97928 272852 97980
rect 282920 97928 282972 97980
rect 283472 97928 283524 97980
rect 284300 97928 284352 97980
rect 284944 97928 284996 97980
rect 285680 97928 285732 97980
rect 286416 97928 286468 97980
rect 287152 97928 287204 97980
rect 288348 97928 288400 97980
rect 291200 97928 291252 97980
rect 291752 97928 291804 97980
rect 292580 97928 292632 97980
rect 293224 97928 293276 97980
rect 293960 97928 294012 97980
rect 294696 97928 294748 97980
rect 295340 97928 295392 97980
rect 296168 97928 296220 97980
rect 299480 97928 299532 97980
rect 300032 97928 300084 97980
rect 300860 97928 300912 97980
rect 301504 97928 301556 97980
rect 302240 97928 302292 97980
rect 302976 97928 303028 97980
rect 303620 97928 303672 97980
rect 304448 97928 304500 97980
rect 307760 97928 307812 97980
rect 308772 97928 308824 97980
rect 309140 97928 309192 97980
rect 310244 97928 310296 97980
rect 310520 97928 310572 97980
rect 311716 97928 311768 97980
rect 311900 97928 311952 97980
rect 313188 97928 313240 97980
rect 317420 97928 317472 97980
rect 318064 97928 318116 97980
rect 318800 97928 318852 97980
rect 319536 97928 319588 97980
rect 320180 97928 320232 97980
rect 321008 97928 321060 97980
rect 321560 97928 321612 97980
rect 322480 97928 322532 97980
rect 324320 97928 324372 97980
rect 324872 97928 324924 97980
rect 327080 97928 327132 97980
rect 327816 97928 327868 97980
rect 328460 97928 328512 97980
rect 329288 97928 329340 97980
rect 92664 97860 92716 97912
rect 93124 97860 93176 97912
rect 98000 97860 98052 97912
rect 98460 97860 98512 97912
rect 116032 97860 116084 97912
rect 116952 97860 117004 97912
rect 136824 97860 136876 97912
rect 137928 97860 137980 97912
rect 140872 97860 140924 97912
rect 141332 97860 141384 97912
rect 176844 97860 176896 97912
rect 177856 97860 177908 97912
rect 197452 97860 197504 97912
rect 198280 97860 198332 97912
rect 198924 97860 198976 97912
rect 199752 97860 199804 97912
rect 215484 97860 215536 97912
rect 216312 97860 216364 97912
rect 216772 97860 216824 97912
rect 217784 97860 217836 97912
rect 218152 97860 218204 97912
rect 219256 97860 219308 97912
rect 220912 97860 220964 97912
rect 222108 97860 222160 97912
rect 229284 97860 229336 97912
rect 230388 97860 230440 97912
rect 231860 97860 231912 97912
rect 232044 97860 232096 97912
rect 237472 97860 237524 97912
rect 238668 97860 238720 97912
rect 249892 97860 249944 97912
rect 250904 97860 250956 97912
rect 256700 97860 256752 97912
rect 257712 97860 257764 97912
rect 289912 97860 289964 97912
rect 290832 97860 290884 97912
rect 291292 97860 291344 97912
rect 292304 97860 292356 97912
rect 298100 97860 298152 97912
rect 298560 97860 298612 97912
rect 306380 97860 306432 97912
rect 307392 97860 307444 97912
rect 323032 97860 323084 97912
rect 323952 97860 324004 97912
rect 324412 97860 324464 97912
rect 325332 97860 325384 97912
rect 106372 97792 106424 97844
rect 107292 97792 107344 97844
rect 107752 97792 107804 97844
rect 108672 97792 108724 97844
rect 180800 97792 180852 97844
rect 181260 97792 181312 97844
rect 182272 97792 182324 97844
rect 182732 97792 182784 97844
rect 183652 97792 183704 97844
rect 184204 97792 184256 97844
rect 197360 97792 197412 97844
rect 197820 97792 197872 97844
rect 200212 97792 200264 97844
rect 201224 97792 201276 97844
rect 240140 97792 240192 97844
rect 240692 97792 240744 97844
rect 243084 97792 243136 97844
rect 244096 97792 244148 97844
rect 281632 97792 281684 97844
rect 282552 97792 282604 97844
rect 283012 97792 283064 97844
rect 284024 97792 284076 97844
rect 289820 97792 289872 97844
rect 290280 97792 290332 97844
rect 322940 97792 322992 97844
rect 323400 97792 323452 97844
rect 128544 97724 128596 97776
rect 129648 97724 129700 97776
rect 219624 97724 219676 97776
rect 220728 97724 220780 97776
rect 231860 97724 231912 97776
rect 232872 97724 232924 97776
rect 245844 97724 245896 97776
rect 246948 97724 247000 97776
rect 281540 97724 281592 97776
rect 282000 97724 282052 97776
rect 106280 96976 106332 97028
rect 106556 96976 106608 97028
rect 147772 94528 147824 94580
rect 148140 94528 148192 94580
rect 150532 94528 150584 94580
rect 151544 94528 151596 94580
rect 154580 94528 154632 94580
rect 155408 94528 155460 94580
rect 155960 94528 156012 94580
rect 156420 94528 156472 94580
rect 3148 85484 3200 85536
rect 90732 85484 90784 85536
rect 577596 73108 577648 73160
rect 579712 73108 579764 73160
rect 3424 71680 3476 71732
rect 90640 71680 90692 71732
rect 92020 60664 92072 60716
rect 580172 60664 580224 60716
rect 3056 59304 3108 59356
rect 90456 59304 90508 59356
rect 3424 45500 3476 45552
rect 90548 45500 90600 45552
rect 3148 33056 3200 33108
rect 90364 33056 90416 33108
rect 577504 33056 577556 33108
rect 579620 33056 579672 33108
rect 254124 23128 254176 23180
rect 393320 23128 393372 23180
rect 256884 23060 256936 23112
rect 400220 23060 400272 23112
rect 259644 22992 259696 23044
rect 407120 22992 407172 23044
rect 262404 22924 262456 22976
rect 415400 22924 415452 22976
rect 265164 22856 265216 22908
rect 422300 22856 422352 22908
rect 267924 22788 267976 22840
rect 429200 22788 429252 22840
rect 270684 22720 270736 22772
rect 436100 22720 436152 22772
rect 240324 22040 240376 22092
rect 361580 22040 361632 22092
rect 241704 21972 241756 22024
rect 365720 21972 365772 22024
rect 243084 21904 243136 21956
rect 368480 21904 368532 21956
rect 244464 21836 244516 21888
rect 372620 21836 372672 21888
rect 245844 21768 245896 21820
rect 375380 21768 375432 21820
rect 248604 21700 248656 21752
rect 379520 21700 379572 21752
rect 249984 21632 250036 21684
rect 382280 21632 382332 21684
rect 251364 21564 251416 21616
rect 386420 21564 386472 21616
rect 309324 21496 309376 21548
rect 528560 21496 528612 21548
rect 310704 21428 310756 21480
rect 531320 21428 531372 21480
rect 312084 21360 312136 21412
rect 535460 21360 535512 21412
rect 238852 21292 238904 21344
rect 357440 21292 357492 21344
rect 237564 21224 237616 21276
rect 354680 21224 354732 21276
rect 236184 21156 236236 21208
rect 350540 21156 350592 21208
rect 92112 20612 92164 20664
rect 579988 20612 580040 20664
rect 252652 20544 252704 20596
rect 391940 20544 391992 20596
rect 254032 20476 254084 20528
rect 396080 20476 396132 20528
rect 256792 20408 256844 20460
rect 398840 20408 398892 20460
rect 258172 20340 258224 20392
rect 402980 20340 403032 20392
rect 278964 20272 279016 20324
rect 456892 20272 456944 20324
rect 281724 20204 281776 20256
rect 459560 20204 459612 20256
rect 283104 20136 283156 20188
rect 463700 20136 463752 20188
rect 284484 20068 284536 20120
rect 466460 20068 466512 20120
rect 285864 20000 285916 20052
rect 470600 20000 470652 20052
rect 307944 19932 307996 19984
rect 524420 19932 524472 19984
rect 251272 19864 251324 19916
rect 389180 19864 389232 19916
rect 234804 19796 234856 19848
rect 347780 19796 347832 19848
rect 232044 19728 232096 19780
rect 339500 19728 339552 19780
rect 267832 19252 267884 19304
rect 426440 19252 426492 19304
rect 269212 19184 269264 19236
rect 430580 19184 430632 19236
rect 270592 19116 270644 19168
rect 433340 19116 433392 19168
rect 271972 19048 272024 19100
rect 437480 19048 437532 19100
rect 298284 18980 298336 19032
rect 502340 18980 502392 19032
rect 299664 18912 299716 18964
rect 506480 18912 506532 18964
rect 301044 18844 301096 18896
rect 509240 18844 509292 18896
rect 302424 18776 302476 18828
rect 513380 18776 513432 18828
rect 303804 18708 303856 18760
rect 516140 18708 516192 18760
rect 325884 18640 325936 18692
rect 569960 18640 570012 18692
rect 327264 18572 327316 18624
rect 572720 18572 572772 18624
rect 266452 18504 266504 18556
rect 423680 18504 423732 18556
rect 229284 18436 229336 18488
rect 335360 18436 335412 18488
rect 227904 18368 227956 18420
rect 332600 18368 332652 18420
rect 242992 17892 243044 17944
rect 365812 17892 365864 17944
rect 244372 17824 244424 17876
rect 369860 17824 369912 17876
rect 290004 17756 290056 17808
rect 480260 17756 480312 17808
rect 291384 17688 291436 17740
rect 483020 17688 483072 17740
rect 292764 17620 292816 17672
rect 487160 17620 487212 17672
rect 294144 17552 294196 17604
rect 489920 17552 489972 17604
rect 295524 17484 295576 17536
rect 494060 17484 494112 17536
rect 317604 17416 317656 17468
rect 547880 17416 547932 17468
rect 318984 17348 319036 17400
rect 550640 17348 550692 17400
rect 320364 17280 320416 17332
rect 554780 17280 554832 17332
rect 321652 17212 321704 17264
rect 557540 17212 557592 17264
rect 241612 17144 241664 17196
rect 362960 17144 363012 17196
rect 240232 17076 240284 17128
rect 358820 17076 358872 17128
rect 237472 17008 237524 17060
rect 356060 17008 356112 17060
rect 233424 16532 233476 16584
rect 344560 16532 344612 16584
rect 313372 16464 313424 16516
rect 539600 16464 539652 16516
rect 314844 16396 314896 16448
rect 542728 16396 542780 16448
rect 316224 16328 316276 16380
rect 546500 16328 546552 16380
rect 317512 16260 317564 16312
rect 550272 16260 550324 16312
rect 318892 16192 318944 16244
rect 553768 16192 553820 16244
rect 323124 16124 323176 16176
rect 560392 16124 560444 16176
rect 324504 16056 324556 16108
rect 564440 16056 564492 16108
rect 325792 15988 325844 16040
rect 567568 15988 567620 16040
rect 327172 15920 327224 15972
rect 571340 15920 571392 15972
rect 216864 15852 216916 15904
rect 303896 15852 303948 15904
rect 328552 15852 328604 15904
rect 575112 15852 575164 15904
rect 231952 15784 232004 15836
rect 340972 15784 341024 15836
rect 230572 15716 230624 15768
rect 337016 15716 337068 15768
rect 229192 15648 229244 15700
rect 332692 15648 332744 15700
rect 289912 15104 289964 15156
rect 482376 15104 482428 15156
rect 291292 15036 291344 15088
rect 486424 15036 486476 15088
rect 292672 14968 292724 15020
rect 490012 14968 490064 15020
rect 294052 14900 294104 14952
rect 493048 14900 493100 14952
rect 298192 14832 298244 14884
rect 500592 14832 500644 14884
rect 295432 14764 295484 14816
rect 497096 14764 497148 14816
rect 299572 14696 299624 14748
rect 503720 14696 503772 14748
rect 300952 14628 301004 14680
rect 507216 14628 507268 14680
rect 302332 14560 302384 14612
rect 511264 14560 511316 14612
rect 303712 14492 303764 14544
rect 514760 14492 514812 14544
rect 305092 14424 305144 14476
rect 517888 14424 517940 14476
rect 288532 14356 288584 14408
rect 478144 14356 478196 14408
rect 287244 14288 287296 14340
rect 474096 14288 474148 14340
rect 227812 14220 227864 14272
rect 330392 14220 330444 14272
rect 263600 13744 263652 13796
rect 417424 13744 417476 13796
rect 265072 13676 265124 13728
rect 420920 13676 420972 13728
rect 266360 13608 266412 13660
rect 423772 13608 423824 13660
rect 267740 13540 267792 13592
rect 428464 13540 428516 13592
rect 269120 13472 269172 13524
rect 432052 13472 432104 13524
rect 270500 13404 270552 13456
rect 435088 13404 435140 13456
rect 271880 13336 271932 13388
rect 439136 13336 439188 13388
rect 273444 13268 273496 13320
rect 442632 13268 442684 13320
rect 274824 13200 274876 13252
rect 445760 13200 445812 13252
rect 276204 13132 276256 13184
rect 448520 13132 448572 13184
rect 277584 13064 277636 13116
rect 453304 13064 453356 13116
rect 262312 12996 262364 13048
rect 414296 12996 414348 13048
rect 260932 12928 260984 12980
rect 410800 12928 410852 12980
rect 259552 12860 259604 12912
rect 407212 12860 407264 12912
rect 236092 12384 236144 12436
rect 349160 12384 349212 12436
rect 237380 12316 237432 12368
rect 353576 12316 353628 12368
rect 238760 12248 238812 12300
rect 357532 12248 357584 12300
rect 240140 12180 240192 12232
rect 361120 12180 361172 12232
rect 241520 12112 241572 12164
rect 364616 12112 364668 12164
rect 242900 12044 242952 12096
rect 367744 12044 367796 12096
rect 244280 11976 244332 12028
rect 371240 11976 371292 12028
rect 245752 11908 245804 11960
rect 374000 11908 374052 11960
rect 247132 11840 247184 11892
rect 378416 11840 378468 11892
rect 248512 11772 248564 11824
rect 382372 11772 382424 11824
rect 249892 11704 249944 11756
rect 385960 11704 386012 11756
rect 110420 11636 110472 11688
rect 110604 11636 110656 11688
rect 234712 11636 234764 11688
rect 346952 11636 347004 11688
rect 233332 11568 233384 11620
rect 342904 11568 342956 11620
rect 226524 11500 226576 11552
rect 326344 11500 326396 11552
rect 284300 11432 284352 11484
rect 284484 11432 284536 11484
rect 309232 10956 309284 11008
rect 527824 10956 527876 11008
rect 214104 10888 214156 10940
rect 298192 10888 298244 10940
rect 310612 10888 310664 10940
rect 531412 10888 531464 10940
rect 215484 10820 215536 10872
rect 301504 10820 301556 10872
rect 311992 10820 312044 10872
rect 534448 10820 534500 10872
rect 216772 10752 216824 10804
rect 305552 10752 305604 10804
rect 313280 10752 313332 10804
rect 538220 10752 538272 10804
rect 218244 10684 218296 10736
rect 307944 10684 307996 10736
rect 314752 10684 314804 10736
rect 541992 10684 542044 10736
rect 218152 10616 218204 10668
rect 309048 10616 309100 10668
rect 316132 10616 316184 10668
rect 545488 10616 545540 10668
rect 219532 10548 219584 10600
rect 311440 10548 311492 10600
rect 317420 10548 317472 10600
rect 548616 10548 548668 10600
rect 219624 10480 219676 10532
rect 312176 10480 312228 10532
rect 318800 10480 318852 10532
rect 552664 10480 552716 10532
rect 221004 10412 221056 10464
rect 314752 10412 314804 10464
rect 320180 10412 320232 10464
rect 556252 10412 556304 10464
rect 222200 10344 222252 10396
rect 318064 10344 318116 10396
rect 323032 10344 323084 10396
rect 563060 10344 563112 10396
rect 220912 10276 220964 10328
rect 316224 10276 316276 10328
rect 324412 10276 324464 10328
rect 566832 10276 566884 10328
rect 307852 10208 307904 10260
rect 523776 10208 523828 10260
rect 306472 10140 306524 10192
rect 520280 10140 520332 10192
rect 226432 10072 226484 10124
rect 328736 10072 328788 10124
rect 225144 10004 225196 10056
rect 324412 10004 324464 10056
rect 225052 9936 225104 9988
rect 323032 9936 323084 9988
rect 223580 9868 223632 9920
rect 319720 9868 319772 9920
rect 278872 9596 278924 9648
rect 455696 9596 455748 9648
rect 280252 9528 280304 9580
rect 459192 9528 459244 9580
rect 281632 9460 281684 9512
rect 462780 9460 462832 9512
rect 283012 9392 283064 9444
rect 466276 9392 466328 9444
rect 85672 9324 85724 9376
rect 127164 9324 127216 9376
rect 203156 9324 203208 9376
rect 270040 9324 270092 9376
rect 285772 9324 285824 9376
rect 473452 9324 473504 9376
rect 45468 9256 45520 9308
rect 110880 9256 110932 9308
rect 204260 9256 204312 9308
rect 273628 9256 273680 9308
rect 287152 9256 287204 9308
rect 476948 9256 477000 9308
rect 41880 9188 41932 9240
rect 109132 9188 109184 9240
rect 205640 9188 205692 9240
rect 277124 9188 277176 9240
rect 289820 9188 289872 9240
rect 481732 9188 481784 9240
rect 38384 9120 38436 9172
rect 107844 9120 107896 9172
rect 207112 9120 207164 9172
rect 280712 9120 280764 9172
rect 291200 9120 291252 9172
rect 485228 9120 485280 9172
rect 34796 9052 34848 9104
rect 106464 9052 106516 9104
rect 208492 9052 208544 9104
rect 284300 9052 284352 9104
rect 292580 9052 292632 9104
rect 488816 9052 488868 9104
rect 31300 8984 31352 9036
rect 103612 8984 103664 9036
rect 209872 8984 209924 9036
rect 287796 8984 287848 9036
rect 293960 8984 294012 9036
rect 492312 8984 492364 9036
rect 27712 8916 27764 8968
rect 102232 8916 102284 8968
rect 211252 8916 211304 8968
rect 291384 8916 291436 8968
rect 296812 8916 296864 8968
rect 499396 8916 499448 8968
rect 276112 8848 276164 8900
rect 448612 8848 448664 8900
rect 273352 8780 273404 8832
rect 441528 8780 441580 8832
rect 215392 8712 215444 8764
rect 300768 8712 300820 8764
rect 214012 8644 214064 8696
rect 297272 8644 297324 8696
rect 212540 8576 212592 8628
rect 294880 8576 294932 8628
rect 51356 8236 51408 8288
rect 111984 8236 112036 8288
rect 249800 8236 249852 8288
rect 384764 8236 384816 8288
rect 47860 8168 47912 8220
rect 110788 8168 110840 8220
rect 251180 8168 251232 8220
rect 388260 8168 388312 8220
rect 33600 8100 33652 8152
rect 105084 8100 105136 8152
rect 201592 8100 201644 8152
rect 237380 8100 237432 8152
rect 252560 8100 252612 8152
rect 391848 8100 391900 8152
rect 30104 8032 30156 8084
rect 103704 8032 103756 8084
rect 203064 8032 203116 8084
rect 240140 8032 240192 8084
rect 253940 8032 253992 8084
rect 395344 8032 395396 8084
rect 26516 7964 26568 8016
rect 102324 7964 102376 8016
rect 207020 7964 207072 8016
rect 249800 7964 249852 8016
rect 255320 7964 255372 8016
rect 398932 7964 398984 8016
rect 23020 7896 23072 7948
rect 100944 7896 100996 7948
rect 187792 7896 187844 7948
rect 234712 7896 234764 7948
rect 256700 7896 256752 7948
rect 402520 7896 402572 7948
rect 18236 7828 18288 7880
rect 99472 7828 99524 7880
rect 193496 7828 193548 7880
rect 248788 7828 248840 7880
rect 258080 7828 258132 7880
rect 406016 7828 406068 7880
rect 7656 7760 7708 7812
rect 94044 7760 94096 7812
rect 194692 7760 194744 7812
rect 251180 7760 251232 7812
rect 259460 7760 259512 7812
rect 409604 7760 409656 7812
rect 2872 7692 2924 7744
rect 92664 7692 92716 7744
rect 201500 7692 201552 7744
rect 258080 7692 258132 7744
rect 260840 7692 260892 7744
rect 413100 7692 413152 7744
rect 572 7624 624 7676
rect 91100 7624 91152 7676
rect 91560 7624 91612 7676
rect 128544 7624 128596 7676
rect 197544 7624 197596 7676
rect 255872 7624 255924 7676
rect 262220 7624 262272 7676
rect 416688 7624 416740 7676
rect 1676 7556 1728 7608
rect 92756 7556 92808 7608
rect 98644 7556 98696 7608
rect 132592 7556 132644 7608
rect 198924 7556 198976 7608
rect 261760 7556 261812 7608
rect 264980 7556 265032 7608
rect 420184 7556 420236 7608
rect 54944 7488 54996 7540
rect 114652 7488 114704 7540
rect 248420 7488 248472 7540
rect 381176 7488 381228 7540
rect 84476 7420 84528 7472
rect 125784 7420 125836 7472
rect 247040 7420 247092 7472
rect 377680 7420 377732 7472
rect 87972 7352 88024 7404
rect 127072 7352 127124 7404
rect 245660 7352 245712 7404
rect 374092 7352 374144 7404
rect 200212 7284 200264 7336
rect 265348 7284 265400 7336
rect 200304 7216 200356 7268
rect 262956 7216 263008 7268
rect 73804 6808 73856 6860
rect 121644 6808 121696 6860
rect 185032 6808 185084 6860
rect 227536 6808 227588 6860
rect 231860 6808 231912 6860
rect 342168 6808 342220 6860
rect 70308 6740 70360 6792
rect 120172 6740 120224 6792
rect 185124 6740 185176 6792
rect 226432 6740 226484 6792
rect 233240 6740 233292 6792
rect 345756 6740 345808 6792
rect 66720 6672 66772 6724
rect 118884 6672 118936 6724
rect 186504 6672 186556 6724
rect 229836 6672 229888 6724
rect 234620 6672 234672 6724
rect 349252 6672 349304 6724
rect 63224 6604 63276 6656
rect 117504 6604 117556 6656
rect 187700 6604 187752 6656
rect 233424 6604 233476 6656
rect 274732 6604 274784 6656
rect 445024 6604 445076 6656
rect 59636 6536 59688 6588
rect 116216 6536 116268 6588
rect 189356 6536 189408 6588
rect 237012 6536 237064 6588
rect 277492 6536 277544 6588
rect 452108 6536 452160 6588
rect 56048 6468 56100 6520
rect 114744 6468 114796 6520
rect 190644 6468 190696 6520
rect 240508 6468 240560 6520
rect 284392 6468 284444 6520
rect 469864 6468 469916 6520
rect 52552 6400 52604 6452
rect 113272 6400 113324 6452
rect 193404 6400 193456 6452
rect 247592 6400 247644 6452
rect 322940 6400 322992 6452
rect 562048 6400 562100 6452
rect 48964 6332 49016 6384
rect 111892 6332 111944 6384
rect 196072 6332 196124 6384
rect 254676 6332 254728 6384
rect 324320 6332 324372 6384
rect 565636 6332 565688 6384
rect 44272 6264 44324 6316
rect 109224 6264 109276 6316
rect 197452 6264 197504 6316
rect 258264 6264 258316 6316
rect 325700 6264 325752 6316
rect 569132 6264 569184 6316
rect 40684 6196 40736 6248
rect 107752 6196 107804 6248
rect 192024 6196 192076 6248
rect 244096 6196 244148 6248
rect 246304 6196 246356 6248
rect 322112 6196 322164 6248
rect 327080 6196 327132 6248
rect 572720 6196 572772 6248
rect 37188 6128 37240 6180
rect 106372 6128 106424 6180
rect 183836 6128 183888 6180
rect 222752 6128 222804 6180
rect 224960 6128 225012 6180
rect 324320 6128 324372 6180
rect 328460 6128 328512 6180
rect 576308 6128 576360 6180
rect 77392 6060 77444 6112
rect 123024 6060 123076 6112
rect 180892 6060 180944 6112
rect 215668 6060 215720 6112
rect 230480 6060 230532 6112
rect 338672 6060 338724 6112
rect 80888 5992 80940 6044
rect 124404 5992 124456 6044
rect 186412 5992 186464 6044
rect 218060 5992 218112 6044
rect 229100 5992 229152 6044
rect 335084 5992 335136 6044
rect 95148 5924 95200 5976
rect 131304 5924 131356 5976
rect 185216 5924 185268 5976
rect 216772 5924 216824 5976
rect 227720 5924 227772 5976
rect 331588 5924 331640 5976
rect 333244 5924 333296 5976
rect 418988 5924 419040 5976
rect 226340 5856 226392 5908
rect 328000 5856 328052 5908
rect 243636 5788 243688 5840
rect 293684 5788 293736 5840
rect 238024 5720 238076 5772
rect 283104 5720 283156 5772
rect 79692 5448 79744 5500
rect 124312 5448 124364 5500
rect 197360 5448 197412 5500
rect 257068 5448 257120 5500
rect 257344 5448 257396 5500
rect 290188 5448 290240 5500
rect 299480 5448 299532 5500
rect 505376 5448 505428 5500
rect 76196 5380 76248 5432
rect 122932 5380 122984 5432
rect 168472 5380 168524 5432
rect 187332 5380 187384 5432
rect 198832 5380 198884 5432
rect 260656 5380 260708 5432
rect 300860 5380 300912 5432
rect 508872 5380 508924 5432
rect 72608 5312 72660 5364
rect 121552 5312 121604 5364
rect 169944 5312 169996 5364
rect 190828 5312 190880 5364
rect 202972 5312 203024 5364
rect 271236 5312 271288 5364
rect 302240 5312 302292 5364
rect 512460 5312 512512 5364
rect 69112 5244 69164 5296
rect 120264 5244 120316 5296
rect 171140 5244 171192 5296
rect 194416 5244 194468 5296
rect 208400 5244 208452 5296
rect 285404 5244 285456 5296
rect 303620 5244 303672 5296
rect 515956 5244 516008 5296
rect 62028 5176 62080 5228
rect 117412 5176 117464 5228
rect 172612 5176 172664 5228
rect 197912 5176 197964 5228
rect 209780 5176 209832 5228
rect 288992 5176 289044 5228
rect 305000 5176 305052 5228
rect 519544 5176 519596 5228
rect 58440 5108 58492 5160
rect 116124 5108 116176 5160
rect 117228 5108 117280 5160
rect 136824 5108 136876 5160
rect 173992 5108 174044 5160
rect 201500 5108 201552 5160
rect 213920 5108 213972 5160
rect 296076 5108 296128 5160
rect 306380 5108 306432 5160
rect 523040 5108 523092 5160
rect 21824 5040 21876 5092
rect 100852 5040 100904 5092
rect 118608 5040 118660 5092
rect 139492 5040 139544 5092
rect 175372 5040 175424 5092
rect 205088 5040 205140 5092
rect 211160 5040 211212 5092
rect 292580 5040 292632 5092
rect 307760 5040 307812 5092
rect 526628 5040 526680 5092
rect 17040 4972 17092 5024
rect 98184 4972 98236 5024
rect 104532 4972 104584 5024
rect 133972 4972 134024 5024
rect 176844 4972 176896 5024
rect 208584 4972 208636 5024
rect 215300 4972 215352 5024
rect 299664 4972 299716 5024
rect 309140 4972 309192 5024
rect 530124 4972 530176 5024
rect 12348 4904 12400 4956
rect 96620 4904 96672 4956
rect 101036 4904 101088 4956
rect 132684 4904 132736 4956
rect 178224 4904 178276 4956
rect 209780 4904 209832 4956
rect 216680 4904 216732 4956
rect 303160 4904 303212 4956
rect 310520 4904 310572 4956
rect 533712 4904 533764 4956
rect 8760 4836 8812 4888
rect 95332 4836 95384 4888
rect 97448 4836 97500 4888
rect 131212 4836 131264 4888
rect 178132 4836 178184 4888
rect 212172 4836 212224 4888
rect 218152 4836 218204 4888
rect 306748 4836 306800 4888
rect 314660 4836 314712 4888
rect 540796 4836 540848 4888
rect 4068 4768 4120 4820
rect 92572 4768 92624 4820
rect 93952 4768 94004 4820
rect 129832 4768 129884 4820
rect 180800 4768 180852 4820
rect 216864 4768 216916 4820
rect 220820 4768 220872 4820
rect 313832 4768 313884 4820
rect 316040 4768 316092 4820
rect 544384 4768 544436 4820
rect 83280 4700 83332 4752
rect 125692 4700 125744 4752
rect 193312 4700 193364 4752
rect 246396 4700 246448 4752
rect 257436 4700 257488 4752
rect 286600 4700 286652 4752
rect 298100 4700 298152 4752
rect 501788 4700 501840 4752
rect 86868 4632 86920 4684
rect 126980 4632 127032 4684
rect 191932 4632 191984 4684
rect 242900 4632 242952 4684
rect 296720 4632 296772 4684
rect 498200 4632 498252 4684
rect 90364 4564 90416 4616
rect 128452 4564 128504 4616
rect 183652 4564 183704 4616
rect 221740 4564 221792 4616
rect 243544 4564 243596 4616
rect 320916 4564 320968 4616
rect 115204 4496 115256 4548
rect 135352 4496 135404 4548
rect 182364 4496 182416 4548
rect 219256 4496 219308 4548
rect 242164 4496 242216 4548
rect 317328 4496 317380 4548
rect 190552 4428 190604 4480
rect 222476 4428 222528 4480
rect 243452 4156 243504 4208
rect 67916 4088 67968 4140
rect 118700 4088 118752 4140
rect 130568 4088 130620 4140
rect 144920 4088 144972 4140
rect 158996 4088 159048 4140
rect 163688 4088 163740 4140
rect 172520 4088 172572 4140
rect 195612 4088 195664 4140
rect 199384 4088 199436 4140
rect 202696 4088 202748 4140
rect 220084 4088 220136 4140
rect 220544 4088 220596 4140
rect 232504 4088 232556 4140
rect 243636 4088 243688 4140
rect 268844 4088 268896 4140
rect 277400 4088 277452 4140
rect 450912 4088 450964 4140
rect 60832 4020 60884 4072
rect 116032 4020 116084 4072
rect 129372 4020 129424 4072
rect 145012 4020 145064 4072
rect 160100 4020 160152 4072
rect 168380 4020 168432 4072
rect 173900 4020 173952 4072
rect 199108 4020 199160 4072
rect 215944 4020 215996 4072
rect 225144 4020 225196 4072
rect 226984 4020 227036 4072
rect 264152 4020 264204 4072
rect 278780 4020 278832 4072
rect 454500 4020 454552 4072
rect 53748 3952 53800 4004
rect 113180 3952 113232 4004
rect 126980 3952 127032 4004
rect 143632 3952 143684 4004
rect 161572 3952 161624 4004
rect 171968 3952 172020 4004
rect 176752 3952 176804 4004
rect 206192 3952 206244 4004
rect 216772 3952 216824 4004
rect 228732 3952 228784 4004
rect 229744 3952 229796 4004
rect 267740 3952 267792 4004
rect 280160 3952 280212 4004
rect 458088 3952 458140 4004
rect 46664 3884 46716 3936
rect 110420 3884 110472 3936
rect 125876 3884 125928 3936
rect 143724 3884 143776 3936
rect 162860 3884 162912 3936
rect 173164 3884 173216 3936
rect 179420 3884 179472 3936
rect 213368 3884 213420 3936
rect 218060 3884 218112 3936
rect 232228 3884 232280 3936
rect 235264 3884 235316 3936
rect 39580 3816 39632 3868
rect 107660 3816 107712 3868
rect 123484 3816 123536 3868
rect 142252 3816 142304 3868
rect 162952 3816 163004 3868
rect 174268 3816 174320 3868
rect 182272 3816 182324 3868
rect 220452 3816 220504 3868
rect 220544 3816 220596 3868
rect 235816 3816 235868 3868
rect 237380 3816 237432 3868
rect 243452 3816 243504 3868
rect 243636 3884 243688 3936
rect 274824 3884 274876 3936
rect 281540 3884 281592 3936
rect 461584 3884 461636 3936
rect 278320 3816 278372 3868
rect 282920 3816 282972 3868
rect 465172 3816 465224 3868
rect 32404 3748 32456 3800
rect 104992 3748 105044 3800
rect 121092 3748 121144 3800
rect 140780 3748 140832 3800
rect 142436 3748 142488 3800
rect 150624 3748 150676 3800
rect 164240 3748 164292 3800
rect 176660 3748 176712 3800
rect 186320 3748 186372 3800
rect 231032 3748 231084 3800
rect 233884 3748 233936 3800
rect 281908 3748 281960 3800
rect 284484 3748 284536 3800
rect 468668 3748 468720 3800
rect 24216 3680 24268 3732
rect 100760 3680 100812 3732
rect 111616 3680 111668 3732
rect 117228 3680 117280 3732
rect 119896 3680 119948 3732
rect 140872 3680 140924 3732
rect 15936 3612 15988 3664
rect 98000 3612 98052 3664
rect 118792 3612 118844 3664
rect 140964 3612 141016 3664
rect 141240 3612 141292 3664
rect 149152 3680 149204 3732
rect 157524 3680 157576 3732
rect 161296 3680 161348 3732
rect 165712 3680 165764 3732
rect 180248 3680 180300 3732
rect 189172 3680 189224 3732
rect 238116 3680 238168 3732
rect 240140 3680 240192 3732
rect 272432 3680 272484 3732
rect 285680 3680 285732 3732
rect 472256 3680 472308 3732
rect 11152 3544 11204 3596
rect 95424 3544 95476 3596
rect 102232 3544 102284 3596
rect 108304 3544 108356 3596
rect 114008 3544 114060 3596
rect 138112 3544 138164 3596
rect 14740 3476 14792 3528
rect 98092 3476 98144 3528
rect 103336 3476 103388 3528
rect 134064 3476 134116 3528
rect 135260 3476 135312 3528
rect 147864 3612 147916 3664
rect 157432 3612 157484 3664
rect 160100 3612 160152 3664
rect 165620 3612 165672 3664
rect 181444 3612 181496 3664
rect 190460 3612 190512 3664
rect 241704 3612 241756 3664
rect 249800 3612 249852 3664
rect 279516 3612 279568 3664
rect 287060 3612 287112 3664
rect 475752 3612 475804 3664
rect 146484 3544 146536 3596
rect 158812 3544 158864 3596
rect 167000 3544 167052 3596
rect 184940 3544 184992 3596
rect 191840 3544 191892 3596
rect 245200 3544 245252 3596
rect 247684 3544 247736 3596
rect 276020 3544 276072 3596
rect 331220 3544 331272 3596
rect 582196 3544 582248 3596
rect 6460 3408 6512 3460
rect 93860 3408 93912 3460
rect 96252 3408 96304 3460
rect 131120 3408 131172 3460
rect 132960 3408 133012 3460
rect 153016 3476 153068 3528
rect 154672 3476 154724 3528
rect 155960 3476 156012 3528
rect 156236 3476 156288 3528
rect 164516 3476 164568 3528
rect 164884 3476 164936 3528
rect 166080 3476 166132 3528
rect 168472 3476 168524 3528
rect 188528 3476 188580 3528
rect 194600 3476 194652 3528
rect 252376 3476 252428 3528
rect 258080 3476 258132 3528
rect 266544 3476 266596 3528
rect 288440 3476 288492 3528
rect 479340 3476 479392 3528
rect 489920 3476 489972 3528
rect 490748 3476 490800 3528
rect 531320 3476 531372 3528
rect 532148 3476 532200 3528
rect 556160 3476 556212 3528
rect 556988 3476 557040 3528
rect 160192 3408 160244 3460
rect 167184 3408 167236 3460
rect 169852 3408 169904 3460
rect 192024 3408 192076 3460
rect 198740 3408 198792 3460
rect 259460 3408 259512 3460
rect 324412 3408 324464 3460
rect 325608 3408 325660 3460
rect 332692 3408 332744 3460
rect 333888 3408 333940 3460
rect 333980 3408 334032 3460
rect 581000 3408 581052 3460
rect 19340 3340 19392 3392
rect 20260 3340 20312 3392
rect 75000 3340 75052 3392
rect 122840 3340 122892 3392
rect 131764 3340 131816 3392
rect 145104 3340 145156 3392
rect 161664 3340 161716 3392
rect 169576 3340 169628 3392
rect 206284 3340 206336 3392
rect 207388 3340 207440 3392
rect 210424 3340 210476 3392
rect 214472 3340 214524 3392
rect 225604 3340 225656 3392
rect 253480 3340 253532 3392
rect 276112 3340 276164 3392
rect 447416 3340 447468 3392
rect 448520 3340 448572 3392
rect 449808 3340 449860 3392
rect 82084 3272 82136 3324
rect 125600 3272 125652 3324
rect 136456 3272 136508 3324
rect 147772 3272 147824 3324
rect 224224 3272 224276 3324
rect 249984 3272 250036 3324
rect 274640 3272 274692 3324
rect 443828 3272 443880 3324
rect 89168 3204 89220 3256
rect 128360 3204 128412 3256
rect 134156 3204 134208 3256
rect 146392 3204 146444 3256
rect 222476 3204 222528 3256
rect 239312 3204 239364 3256
rect 273260 3204 273312 3256
rect 440332 3204 440384 3256
rect 209044 3136 209096 3188
rect 210976 3136 211028 3188
rect 211804 3136 211856 3188
rect 218060 3136 218112 3188
rect 329840 3136 329892 3188
rect 333980 3136 334032 3188
rect 349160 3136 349212 3188
rect 350448 3136 350500 3188
rect 357440 3136 357492 3188
rect 358728 3136 358780 3188
rect 365812 3136 365864 3188
rect 367008 3136 367060 3188
rect 374000 3136 374052 3188
rect 375288 3136 375340 3188
rect 382280 3136 382332 3188
rect 383568 3136 383620 3188
rect 398840 3136 398892 3188
rect 400128 3136 400180 3188
rect 407120 3136 407172 3188
rect 408408 3136 408460 3188
rect 423772 3136 423824 3188
rect 424968 3136 425020 3188
rect 431960 3136 432012 3188
rect 433248 3136 433300 3188
rect 145932 3068 145984 3120
rect 151912 3068 151964 3120
rect 128176 3000 128228 3052
rect 129004 3000 129056 3052
rect 144736 3000 144788 3052
rect 150532 3000 150584 3052
rect 213184 3000 213236 3052
rect 221556 3000 221608 3052
rect 149520 2932 149572 2984
rect 153384 2932 153436 2984
rect 108120 2796 108172 2848
rect 115204 2796 115256 2848
rect 115296 2796 115348 2848
rect 118608 2796 118660 2848
rect 221740 2796 221792 2848
rect 223948 2796 224000 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700466 8156 703520
rect 24320 700534 24348 703520
rect 24308 700528 24360 700534
rect 24308 700470 24360 700476
rect 8116 700460 8168 700466
rect 8116 700402 8168 700408
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683262 3464 684247
rect 3424 683256 3476 683262
rect 3424 683198 3476 683204
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3436 670818 3464 671191
rect 3424 670812 3476 670818
rect 3424 670754 3476 670760
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 422346 3464 423535
rect 3424 422340 3476 422346
rect 3424 422282 3476 422288
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 409902 3188 410479
rect 3148 409896 3200 409902
rect 3148 409838 3200 409844
rect 3424 397520 3476 397526
rect 3422 397488 3424 397497
rect 3476 397488 3478 397497
rect 3422 397423 3478 397432
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 371278 3464 371311
rect 3424 371272 3476 371278
rect 3424 371214 3476 371220
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 40052 346050 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 700738 73016 703520
rect 89180 700806 89208 703520
rect 89168 700800 89220 700806
rect 89168 700742 89220 700748
rect 72976 700732 73028 700738
rect 72976 700674 73028 700680
rect 104912 346186 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 137848 701010 137876 703520
rect 137836 701004 137888 701010
rect 137836 700946 137888 700952
rect 154132 700262 154160 703520
rect 170324 702434 170352 703520
rect 169772 702406 170352 702434
rect 154120 700256 154172 700262
rect 154120 700198 154172 700204
rect 168380 563100 168432 563106
rect 168380 563042 168432 563048
rect 164240 536852 164292 536858
rect 164240 536794 164292 536800
rect 161480 510672 161532 510678
rect 161480 510614 161532 510620
rect 157340 484424 157392 484430
rect 157340 484366 157392 484372
rect 155960 456816 156012 456822
rect 155960 456758 156012 456764
rect 151820 430636 151872 430642
rect 151820 430578 151872 430584
rect 149060 404388 149112 404394
rect 149060 404330 149112 404336
rect 144920 378208 144972 378214
rect 144920 378150 144972 378156
rect 144932 364334 144960 378150
rect 147680 364404 147732 364410
rect 147680 364346 147732 364352
rect 144932 364306 145328 364334
rect 143540 351960 143592 351966
rect 143540 351902 143592 351908
rect 109408 347812 109460 347818
rect 109408 347754 109460 347760
rect 104900 346180 104952 346186
rect 104900 346122 104952 346128
rect 40040 346044 40092 346050
rect 40040 345986 40092 345992
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 99286 344720 99342 344729
rect 99286 344655 99342 344664
rect 90640 344276 90692 344282
rect 90640 344218 90692 344224
rect 3516 344208 3568 344214
rect 3516 344150 3568 344156
rect 3424 344004 3476 344010
rect 3424 343946 3476 343952
rect 3240 341420 3292 341426
rect 3240 341362 3292 341368
rect 3252 319297 3280 341362
rect 3332 341284 3384 341290
rect 3332 341226 3384 341232
rect 3238 319288 3294 319297
rect 3238 319223 3294 319232
rect 3344 306241 3372 341226
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 2780 163804 2832 163810
rect 2780 163746 2832 163752
rect 2792 162897 2820 163746
rect 2778 162888 2834 162897
rect 2778 162823 2834 162832
rect 3436 149841 3464 343946
rect 3528 188873 3556 344150
rect 3608 344140 3660 344146
rect 3608 344082 3660 344088
rect 3620 201929 3648 344082
rect 4896 344072 4948 344078
rect 4896 344014 4948 344020
rect 4804 343936 4856 343942
rect 4804 343878 4856 343884
rect 3976 342644 4028 342650
rect 3976 342586 4028 342592
rect 3700 342576 3752 342582
rect 3700 342518 3752 342524
rect 3712 214985 3740 342518
rect 3792 341216 3844 341222
rect 3792 341158 3844 341164
rect 3804 241097 3832 341158
rect 3884 341148 3936 341154
rect 3884 341090 3936 341096
rect 3896 254153 3924 341090
rect 3988 267209 4016 342586
rect 4068 341352 4120 341358
rect 4068 341294 4120 341300
rect 4080 293185 4108 341294
rect 4066 293176 4122 293185
rect 4066 293111 4122 293120
rect 3974 267200 4030 267209
rect 3974 267135 4030 267144
rect 3882 254144 3938 254153
rect 3882 254079 3938 254088
rect 3790 241088 3846 241097
rect 3790 241023 3846 241032
rect 3698 214976 3754 214985
rect 3698 214911 3754 214920
rect 3606 201920 3662 201929
rect 3606 201855 3662 201864
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 4816 110770 4844 343878
rect 4908 163810 4936 344014
rect 90456 342712 90508 342718
rect 90456 342654 90508 342660
rect 90362 341320 90418 341329
rect 90362 341255 90418 341264
rect 4896 163804 4948 163810
rect 4896 163746 4948 163752
rect 2780 110764 2832 110770
rect 2780 110706 2832 110712
rect 4804 110764 4856 110770
rect 4804 110706 4856 110712
rect 2792 110673 2820 110706
rect 2778 110664 2834 110673
rect 2778 110599 2834 110608
rect 70400 100700 70452 100706
rect 70400 100642 70452 100648
rect 63500 100632 63552 100638
rect 63500 100574 63552 100580
rect 56600 100564 56652 100570
rect 56600 100506 56652 100512
rect 49700 100496 49752 100502
rect 49700 100438 49752 100444
rect 42800 100428 42852 100434
rect 42800 100370 42852 100376
rect 35900 100360 35952 100366
rect 35900 100302 35952 100308
rect 27620 100292 27672 100298
rect 27620 100234 27672 100240
rect 19432 100224 19484 100230
rect 19432 100166 19484 100172
rect 19340 100088 19392 100094
rect 19340 100030 19392 100036
rect 9680 100020 9732 100026
rect 9680 99962 9732 99968
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3148 33108 3200 33114
rect 3148 33050 3200 33056
rect 3160 32473 3188 33050
rect 3146 32464 3202 32473
rect 3146 32399 3202 32408
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 572 7676 624 7682
rect 572 7618 624 7624
rect 584 480 612 7618
rect 1676 7608 1728 7614
rect 1676 7550 1728 7556
rect 1688 480 1716 7550
rect 2884 480 2912 7686
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4080 480 4108 4762
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 5262 3360 5318 3369
rect 5262 3295 5318 3304
rect 5276 480 5304 3295
rect 6472 480 6500 3402
rect 7668 480 7696 7754
rect 8760 4888 8812 4894
rect 8760 4830 8812 4836
rect 8772 480 8800 4830
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 99962
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 13542 6216 13598 6225
rect 13542 6151 13598 6160
rect 12348 4956 12400 4962
rect 12348 4898 12400 4904
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11164 480 11192 3538
rect 12360 480 12388 4898
rect 13556 480 13584 6151
rect 17040 5024 17092 5030
rect 17040 4966 17092 4972
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14752 480 14780 3470
rect 15948 480 15976 3606
rect 17052 480 17080 4966
rect 18248 480 18276 7822
rect 19352 3398 19380 100030
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19444 480 19472 100166
rect 24860 100156 24912 100162
rect 24860 100098 24912 100104
rect 24872 16574 24900 100098
rect 27632 16574 27660 100234
rect 35912 16574 35940 100302
rect 24872 16546 25360 16574
rect 27632 16546 28488 16574
rect 35912 16546 36032 16574
rect 23020 7948 23072 7954
rect 23020 7890 23072 7896
rect 21824 5092 21876 5098
rect 21824 5034 21876 5040
rect 20260 3392 20312 3398
rect 20260 3334 20312 3340
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20272 354 20300 3334
rect 21836 480 21864 5034
rect 23032 480 23060 7890
rect 24216 3732 24268 3738
rect 24216 3674 24268 3680
rect 24228 480 24256 3674
rect 25332 480 25360 16546
rect 27712 8968 27764 8974
rect 27712 8910 27764 8916
rect 26516 8016 26568 8022
rect 26516 7958 26568 7964
rect 26528 480 26556 7958
rect 27724 480 27752 8910
rect 20598 354 20710 480
rect 20272 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 34796 9104 34848 9110
rect 34796 9046 34848 9052
rect 31300 9036 31352 9042
rect 31300 8978 31352 8984
rect 30104 8084 30156 8090
rect 30104 8026 30156 8032
rect 30116 480 30144 8026
rect 31312 480 31340 8978
rect 33600 8152 33652 8158
rect 33600 8094 33652 8100
rect 32404 3800 32456 3806
rect 32404 3742 32456 3748
rect 32416 480 32444 3742
rect 33612 480 33640 8094
rect 34808 480 34836 9046
rect 36004 480 36032 16546
rect 41880 9240 41932 9246
rect 41880 9182 41932 9188
rect 38384 9172 38436 9178
rect 38384 9114 38436 9120
rect 37188 6180 37240 6186
rect 37188 6122 37240 6128
rect 37200 480 37228 6122
rect 38396 480 38424 9114
rect 40684 6248 40736 6254
rect 40684 6190 40736 6196
rect 39580 3868 39632 3874
rect 39580 3810 39632 3816
rect 39592 480 39620 3810
rect 40696 480 40724 6190
rect 41892 480 41920 9182
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 42812 354 42840 100370
rect 49712 16574 49740 100438
rect 56612 16574 56640 100506
rect 63512 16574 63540 100574
rect 70412 16574 70440 100642
rect 77300 99952 77352 99958
rect 77300 99894 77352 99900
rect 77312 16574 77340 99894
rect 90376 33114 90404 341255
rect 90468 59362 90496 342654
rect 90546 341456 90602 341465
rect 90546 341391 90602 341400
rect 90456 59356 90508 59362
rect 90456 59298 90508 59304
rect 90560 45558 90588 341391
rect 90652 71738 90680 344218
rect 92020 343868 92072 343874
rect 92020 343810 92072 343816
rect 90824 342780 90876 342786
rect 90824 342722 90876 342728
rect 90732 341488 90784 341494
rect 90732 341430 90784 341436
rect 90744 85542 90772 341430
rect 90836 97986 90864 342722
rect 90824 97980 90876 97986
rect 90824 97922 90876 97928
rect 91100 97980 91152 97986
rect 91100 97922 91152 97928
rect 90732 85536 90784 85542
rect 90732 85478 90784 85484
rect 90640 71732 90692 71738
rect 90640 71674 90692 71680
rect 90548 45552 90600 45558
rect 90548 45494 90600 45500
rect 90364 33108 90416 33114
rect 90364 33050 90416 33056
rect 49712 16546 50200 16574
rect 56612 16546 56824 16574
rect 63512 16546 64368 16574
rect 70412 16546 71544 16574
rect 77312 16546 78168 16574
rect 45468 9308 45520 9314
rect 45468 9250 45520 9256
rect 44272 6316 44324 6322
rect 44272 6258 44324 6264
rect 44284 480 44312 6258
rect 45480 480 45508 9250
rect 47860 8220 47912 8226
rect 47860 8162 47912 8168
rect 46664 3936 46716 3942
rect 46664 3878 46716 3884
rect 46676 480 46704 3878
rect 47872 480 47900 8162
rect 48964 6384 49016 6390
rect 48964 6326 49016 6332
rect 48976 480 49004 6326
rect 50172 480 50200 16546
rect 51356 8288 51408 8294
rect 51356 8230 51408 8236
rect 51368 480 51396 8230
rect 54944 7540 54996 7546
rect 54944 7482 54996 7488
rect 52552 6452 52604 6458
rect 52552 6394 52604 6400
rect 52564 480 52592 6394
rect 53748 4004 53800 4010
rect 53748 3946 53800 3952
rect 53760 480 53788 3946
rect 54956 480 54984 7482
rect 56048 6520 56100 6526
rect 56048 6462 56100 6468
rect 56060 480 56088 6462
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 63224 6656 63276 6662
rect 63224 6598 63276 6604
rect 59636 6588 59688 6594
rect 59636 6530 59688 6536
rect 58440 5160 58492 5166
rect 58440 5102 58492 5108
rect 58452 480 58480 5102
rect 59648 480 59676 6530
rect 62028 5228 62080 5234
rect 62028 5170 62080 5176
rect 60832 4072 60884 4078
rect 60832 4014 60884 4020
rect 60844 480 60872 4014
rect 62040 480 62068 5170
rect 63236 480 63264 6598
rect 64340 480 64368 16546
rect 70308 6792 70360 6798
rect 70308 6734 70360 6740
rect 66720 6724 66772 6730
rect 66720 6666 66772 6672
rect 65522 4856 65578 4865
rect 65522 4791 65578 4800
rect 65536 480 65564 4791
rect 66732 480 66760 6666
rect 69112 5296 69164 5302
rect 69112 5238 69164 5244
rect 67916 4140 67968 4146
rect 67916 4082 67968 4088
rect 67928 480 67956 4082
rect 69124 480 69152 5238
rect 70320 480 70348 6734
rect 71516 480 71544 16546
rect 73804 6860 73856 6866
rect 73804 6802 73856 6808
rect 72608 5364 72660 5370
rect 72608 5306 72660 5312
rect 72620 480 72648 5306
rect 73816 480 73844 6802
rect 77392 6112 77444 6118
rect 77392 6054 77444 6060
rect 76196 5432 76248 5438
rect 76196 5374 76248 5380
rect 75000 3392 75052 3398
rect 75000 3334 75052 3340
rect 75012 480 75040 3334
rect 76208 480 76236 5374
rect 77404 480 77432 6054
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 85672 9376 85724 9382
rect 85672 9318 85724 9324
rect 84476 7472 84528 7478
rect 84476 7414 84528 7420
rect 80888 6044 80940 6050
rect 80888 5986 80940 5992
rect 79692 5500 79744 5506
rect 79692 5442 79744 5448
rect 79704 480 79732 5442
rect 80900 480 80928 5986
rect 83280 4752 83332 4758
rect 83280 4694 83332 4700
rect 82084 3324 82136 3330
rect 82084 3266 82136 3272
rect 82096 480 82124 3266
rect 83292 480 83320 4694
rect 84488 480 84516 7414
rect 85684 480 85712 9318
rect 91112 7682 91140 97922
rect 92032 60722 92060 343810
rect 92112 343800 92164 343806
rect 92112 343742 92164 343748
rect 97172 343800 97224 343806
rect 97172 343742 97224 343748
rect 92020 60716 92072 60722
rect 92020 60658 92072 60664
rect 92124 20670 92152 343742
rect 95056 343732 95108 343738
rect 95056 343674 95108 343680
rect 93032 343664 93084 343670
rect 93032 343606 93084 343612
rect 93044 341972 93072 343606
rect 95068 341972 95096 343674
rect 97184 341972 97212 343742
rect 99300 341972 99328 344655
rect 103520 343868 103572 343874
rect 103520 343810 103572 343816
rect 105636 343868 105688 343874
rect 105636 343810 105688 343816
rect 101404 343800 101456 343806
rect 101404 343742 101456 343748
rect 101416 341972 101444 343742
rect 103532 341972 103560 343810
rect 105648 341972 105676 343810
rect 109420 341986 109448 347754
rect 141422 344584 141478 344593
rect 141422 344519 141478 344528
rect 135074 344448 135130 344457
rect 126704 344412 126756 344418
rect 135074 344383 135130 344392
rect 126704 344354 126756 344360
rect 114008 344344 114060 344350
rect 114008 344286 114060 344292
rect 111892 342304 111944 342310
rect 111892 342246 111944 342252
rect 109420 341958 109894 341986
rect 111904 341972 111932 342246
rect 114020 341972 114048 344286
rect 116122 344040 116178 344049
rect 116122 343975 116178 343984
rect 116136 341972 116164 343975
rect 124588 342508 124640 342514
rect 124588 342450 124640 342456
rect 122472 342440 122524 342446
rect 122472 342382 122524 342388
rect 118240 342372 118292 342378
rect 118240 342314 118292 342320
rect 118252 341972 118280 342314
rect 122484 341972 122512 342382
rect 124600 341972 124628 342450
rect 126716 341972 126744 344354
rect 132958 344312 133014 344321
rect 132958 344247 133014 344256
rect 128818 344176 128874 344185
rect 128818 344111 128874 344120
rect 128832 341972 128860 344111
rect 132972 341972 133000 344247
rect 135088 341972 135116 344383
rect 141436 341972 141464 344519
rect 143552 341972 143580 351902
rect 145300 341986 145328 364306
rect 147692 341986 147720 364346
rect 149072 364334 149100 404330
rect 149072 364306 149376 364334
rect 149348 341986 149376 364306
rect 151832 341986 151860 430578
rect 153200 418192 153252 418198
rect 153200 418134 153252 418140
rect 153212 364334 153240 418134
rect 153212 364306 153608 364334
rect 153580 341986 153608 364306
rect 155972 341986 156000 456758
rect 157352 364334 157380 484366
rect 160100 470620 160152 470626
rect 160100 470562 160152 470568
rect 157352 364306 157840 364334
rect 157812 341986 157840 364306
rect 160112 341986 160140 470562
rect 161492 364334 161520 510614
rect 161492 364306 162072 364334
rect 162044 341986 162072 364306
rect 164252 341986 164280 536794
rect 165620 524476 165672 524482
rect 165620 524418 165672 524424
rect 165632 364334 165660 524418
rect 165632 364306 166304 364334
rect 166276 341986 166304 364306
rect 168392 341986 168420 563042
rect 169772 346322 169800 702406
rect 201500 700664 201552 700670
rect 201500 700606 201552 700612
rect 197360 700392 197412 700398
rect 197360 700334 197412 700340
rect 191840 700324 191892 700330
rect 191840 700266 191892 700272
rect 183560 696992 183612 696998
rect 183560 696934 183612 696940
rect 180800 670744 180852 670750
rect 180800 670686 180852 670692
rect 176660 643136 176712 643142
rect 176660 643078 176712 643084
rect 173900 616888 173952 616894
rect 173900 616830 173952 616836
rect 169852 590708 169904 590714
rect 169852 590650 169904 590656
rect 169864 364334 169892 590650
rect 172520 576904 172572 576910
rect 172520 576846 172572 576852
rect 169864 364306 170536 364334
rect 169760 346316 169812 346322
rect 169760 346258 169812 346264
rect 170508 341986 170536 364306
rect 172532 341986 172560 576846
rect 173912 364334 173940 616830
rect 176672 364334 176700 643078
rect 178040 630692 178092 630698
rect 178040 630634 178092 630640
rect 178052 364334 178080 630634
rect 180812 364334 180840 670686
rect 173912 364306 174768 364334
rect 176672 364306 176792 364334
rect 178052 364306 179000 364334
rect 180812 364306 181024 364334
rect 174740 341986 174768 364306
rect 176764 341986 176792 364306
rect 178972 341986 179000 364306
rect 180996 341986 181024 364306
rect 145300 341958 145682 341986
rect 147692 341958 147798 341986
rect 149348 341958 149822 341986
rect 151832 341958 151938 341986
rect 153580 341958 154054 341986
rect 155972 341958 156170 341986
rect 157812 341958 158286 341986
rect 160112 341958 160402 341986
rect 162044 341958 162518 341986
rect 164252 341958 164634 341986
rect 166276 341958 166750 341986
rect 168392 341958 168774 341986
rect 170508 341958 170890 341986
rect 172532 341958 173006 341986
rect 174740 341958 175122 341986
rect 176764 341958 177238 341986
rect 178972 341958 179354 341986
rect 180996 341958 181470 341986
rect 183572 341972 183600 696934
rect 184940 683188 184992 683194
rect 184940 683130 184992 683136
rect 184952 364334 184980 683130
rect 184952 364306 185256 364334
rect 185228 341986 185256 364306
rect 189816 345772 189868 345778
rect 189816 345714 189868 345720
rect 187700 345704 187752 345710
rect 187700 345646 187752 345652
rect 185228 341958 185610 341986
rect 187712 341972 187740 345646
rect 189828 341972 189856 345714
rect 191852 341986 191880 700266
rect 197372 364334 197400 700334
rect 201512 364334 201540 700606
rect 202800 700194 202828 703520
rect 208400 700936 208452 700942
rect 208400 700878 208452 700884
rect 204260 700596 204312 700602
rect 204260 700538 204312 700544
rect 202788 700188 202840 700194
rect 202788 700130 202840 700136
rect 197372 364306 197952 364334
rect 201512 364306 202184 364334
rect 196164 345908 196216 345914
rect 196164 345850 196216 345856
rect 194048 345840 194100 345846
rect 194048 345782 194100 345788
rect 191852 341958 191958 341986
rect 194060 341972 194088 345782
rect 196176 341972 196204 345850
rect 197924 341986 197952 364306
rect 200396 345976 200448 345982
rect 200396 345918 200448 345924
rect 197924 341958 198306 341986
rect 200408 341972 200436 345918
rect 202156 341986 202184 364306
rect 204272 341986 204300 700538
rect 206652 346112 206704 346118
rect 206652 346054 206704 346060
rect 202156 341958 202538 341986
rect 204272 341958 204562 341986
rect 206664 341972 206692 346054
rect 208412 341986 208440 700878
rect 209780 700868 209832 700874
rect 209780 700810 209832 700816
rect 209792 364334 209820 700810
rect 215944 700188 215996 700194
rect 215944 700130 215996 700136
rect 216680 700188 216732 700194
rect 216680 700130 216732 700136
rect 209792 364306 210464 364334
rect 210436 341986 210464 364306
rect 215116 346384 215168 346390
rect 215116 346326 215168 346332
rect 213000 346248 213052 346254
rect 213000 346190 213052 346196
rect 208412 341958 208794 341986
rect 210436 341958 210910 341986
rect 213012 341972 213040 346190
rect 215128 341972 215156 346326
rect 215956 344554 215984 700130
rect 216692 364334 216720 700130
rect 218992 700126 219020 703520
rect 227720 701004 227772 701010
rect 227720 700946 227772 700952
rect 218980 700120 219032 700126
rect 218980 700062 219032 700068
rect 222200 700120 222252 700126
rect 222200 700062 222252 700068
rect 222212 364334 222240 700062
rect 216692 364306 216904 364334
rect 222212 364306 223160 364334
rect 215944 344548 215996 344554
rect 215944 344490 215996 344496
rect 216876 341986 216904 364306
rect 219348 345636 219400 345642
rect 219348 345578 219400 345584
rect 216876 341958 217258 341986
rect 219360 341972 219388 345578
rect 220820 345092 220872 345098
rect 220820 345034 220872 345040
rect 220832 344486 220860 345034
rect 221464 344548 221516 344554
rect 221464 344490 221516 344496
rect 220820 344480 220872 344486
rect 220820 344422 220872 344428
rect 221476 341972 221504 344490
rect 223132 341986 223160 364306
rect 225604 346316 225656 346322
rect 225604 346258 225656 346264
rect 223132 341958 223514 341986
rect 225616 341972 225644 346258
rect 227732 341972 227760 700946
rect 233240 700732 233292 700738
rect 233240 700674 233292 700680
rect 229100 700256 229152 700262
rect 229100 700198 229152 700204
rect 229112 364334 229140 700198
rect 233252 364334 233280 700674
rect 229112 364306 229416 364334
rect 233252 364306 233648 364334
rect 229388 341986 229416 364306
rect 231952 346180 232004 346186
rect 231952 346122 232004 346128
rect 229388 341958 229862 341986
rect 231964 341972 231992 346122
rect 233620 341986 233648 364306
rect 234632 345642 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 236000 700800 236052 700806
rect 236000 700742 236052 700748
rect 234620 345636 234672 345642
rect 234620 345578 234672 345584
rect 236012 341986 236040 700742
rect 241520 700528 241572 700534
rect 241520 700470 241572 700476
rect 240140 700460 240192 700466
rect 240140 700402 240192 700408
rect 238300 346044 238352 346050
rect 238300 345986 238352 345992
rect 233620 341958 234094 341986
rect 236012 341958 236210 341986
rect 238312 341972 238340 345986
rect 240152 341986 240180 700402
rect 241532 364334 241560 700470
rect 267660 693530 267688 703520
rect 283852 700194 283880 703520
rect 283840 700188 283892 700194
rect 283840 700130 283892 700136
rect 266360 693524 266412 693530
rect 266360 693466 266412 693472
rect 267648 693524 267700 693530
rect 267648 693466 267700 693472
rect 244280 683256 244332 683262
rect 244280 683198 244332 683204
rect 241532 364306 242112 364334
rect 242084 341986 242112 364306
rect 244292 341986 244320 683198
rect 248420 670812 248472 670818
rect 248420 670754 248472 670760
rect 245660 656940 245712 656946
rect 245660 656882 245712 656888
rect 245672 364334 245700 656882
rect 245672 364306 246344 364334
rect 246316 341986 246344 364306
rect 248432 341986 248460 670754
rect 249800 632120 249852 632126
rect 249800 632062 249852 632068
rect 249812 364334 249840 632062
rect 253940 618316 253992 618322
rect 253940 618258 253992 618264
rect 252560 605872 252612 605878
rect 252560 605814 252612 605820
rect 249812 364306 250576 364334
rect 250548 341986 250576 364306
rect 252572 341986 252600 605814
rect 253952 364334 253980 618258
rect 256700 579692 256752 579698
rect 256700 579634 256752 579640
rect 256712 364334 256740 579634
rect 260840 565888 260892 565894
rect 260840 565830 260892 565836
rect 258080 553444 258132 553450
rect 258080 553386 258132 553392
rect 258092 364334 258120 553386
rect 260852 364334 260880 565830
rect 262220 527196 262272 527202
rect 262220 527138 262272 527144
rect 262232 364334 262260 527138
rect 264980 501016 265032 501022
rect 264980 500958 265032 500964
rect 264992 364334 265020 500958
rect 253952 364306 254808 364334
rect 256712 364306 256832 364334
rect 258092 364306 258856 364334
rect 260852 364306 261064 364334
rect 262232 364306 263088 364334
rect 264992 364306 265296 364334
rect 254780 341986 254808 364306
rect 256804 341986 256832 364306
rect 258828 341986 258856 364306
rect 261036 341986 261064 364306
rect 263060 341986 263088 364306
rect 265268 341986 265296 364306
rect 266372 346390 266400 693466
rect 267740 514820 267792 514826
rect 267740 514762 267792 514768
rect 266360 346384 266412 346390
rect 266360 346326 266412 346332
rect 240152 341958 240442 341986
rect 242084 341958 242466 341986
rect 244292 341958 244582 341986
rect 246316 341958 246698 341986
rect 248432 341958 248814 341986
rect 250548 341958 250930 341986
rect 252572 341958 253046 341986
rect 254780 341958 255162 341986
rect 256804 341958 257278 341986
rect 258828 341958 259302 341986
rect 261036 341958 261418 341986
rect 263060 341958 263534 341986
rect 265268 341958 265650 341986
rect 267752 341972 267780 514762
rect 269120 474768 269172 474774
rect 269120 474710 269172 474716
rect 269132 364334 269160 474710
rect 273260 462392 273312 462398
rect 273260 462334 273312 462340
rect 271880 448588 271932 448594
rect 271880 448530 271932 448536
rect 269132 364306 269528 364334
rect 269500 341986 269528 364306
rect 271892 341986 271920 448530
rect 273272 364334 273300 462334
rect 276020 422340 276072 422346
rect 276020 422282 276072 422288
rect 273272 364306 273760 364334
rect 273732 341986 273760 364306
rect 276032 341986 276060 422282
rect 280160 409896 280212 409902
rect 280160 409838 280212 409844
rect 277400 397520 277452 397526
rect 277400 397462 277452 397468
rect 277412 364334 277440 397462
rect 277412 364306 277808 364334
rect 277780 341986 277808 364306
rect 280172 341986 280200 409838
rect 281540 371272 281592 371278
rect 281540 371214 281592 371220
rect 281552 364334 281580 371214
rect 281552 364306 282040 364334
rect 282012 341986 282040 364306
rect 284944 357468 284996 357474
rect 284944 357410 284996 357416
rect 284956 344486 284984 357410
rect 299492 346254 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 700942 332548 703520
rect 332508 700936 332560 700942
rect 332508 700878 332560 700884
rect 348804 700874 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700868 348844 700874
rect 348792 700810 348844 700816
rect 299480 346248 299532 346254
rect 299480 346190 299532 346196
rect 364352 346118 364380 702406
rect 397472 700670 397500 703520
rect 397460 700664 397512 700670
rect 397460 700606 397512 700612
rect 413664 700602 413692 703520
rect 413652 700596 413704 700602
rect 413652 700538 413704 700544
rect 364340 346112 364392 346118
rect 364340 346054 364392 346060
rect 429212 345982 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 429200 345976 429252 345982
rect 429200 345918 429252 345924
rect 462332 345914 462360 703520
rect 478524 700398 478552 703520
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 462320 345908 462372 345914
rect 462320 345850 462372 345856
rect 494072 345846 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 494060 345840 494112 345846
rect 494060 345782 494112 345788
rect 527192 345778 527220 703520
rect 543476 700330 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 527180 345772 527232 345778
rect 527180 345714 527232 345720
rect 558932 345710 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 577688 347812 577740 347818
rect 577688 347754 577740 347760
rect 558920 345704 558972 345710
rect 558920 345646 558972 345652
rect 284576 344480 284628 344486
rect 284576 344422 284628 344428
rect 284944 344480 284996 344486
rect 284944 344422 284996 344428
rect 286692 344480 286744 344486
rect 286692 344422 286744 344428
rect 269500 341958 269882 341986
rect 271892 341958 271998 341986
rect 273732 341958 274114 341986
rect 276032 341958 276230 341986
rect 277780 341958 278254 341986
rect 280172 341958 280370 341986
rect 282012 341958 282486 341986
rect 284588 341972 284616 344422
rect 286704 341972 286732 344422
rect 331956 344412 332008 344418
rect 331956 344354 332008 344360
rect 331864 344344 331916 344350
rect 331864 344286 331916 344292
rect 320364 344276 320416 344282
rect 320364 344218 320416 344224
rect 303528 344208 303580 344214
rect 303528 344150 303580 344156
rect 295156 342644 295208 342650
rect 295156 342586 295208 342592
rect 295168 341972 295196 342586
rect 301412 342576 301464 342582
rect 301412 342518 301464 342524
rect 301424 341972 301452 342518
rect 303540 341972 303568 344150
rect 305644 344140 305696 344146
rect 305644 344082 305696 344088
rect 305656 341972 305684 344082
rect 307760 344072 307812 344078
rect 307760 344014 307812 344020
rect 307772 341972 307800 344014
rect 311992 344004 312044 344010
rect 311992 343946 312044 343952
rect 309874 343904 309930 343913
rect 309874 343839 309930 343848
rect 309888 341972 309916 343839
rect 312004 341972 312032 343946
rect 314108 343936 314160 343942
rect 314108 343878 314160 343884
rect 314120 341972 314148 343878
rect 318248 342780 318300 342786
rect 318248 342722 318300 342728
rect 318260 341972 318288 342722
rect 320376 341972 320404 344218
rect 324596 342712 324648 342718
rect 324596 342654 324648 342660
rect 324608 341972 324636 342654
rect 135260 341828 135312 341834
rect 135260 341770 135312 341776
rect 164792 341828 164844 341834
rect 164792 341770 164844 341776
rect 135272 341630 135300 341770
rect 135260 341624 135312 341630
rect 108118 341592 108174 341601
rect 107778 341550 108118 341578
rect 120630 341592 120686 341601
rect 120382 341550 120630 341578
rect 108118 341527 108174 341536
rect 135536 341624 135588 341630
rect 135260 341566 135312 341572
rect 135350 341592 135406 341601
rect 120630 341527 120686 341536
rect 135536 341566 135588 341572
rect 139952 341624 140004 341630
rect 139952 341566 140004 341572
rect 164146 341592 164202 341601
rect 135350 341527 135406 341536
rect 135444 341556 135496 341562
rect 135214 341488 135266 341494
rect 130870 341426 131160 341442
rect 135364 341442 135392 341527
rect 135444 341498 135496 341504
rect 135266 341436 135392 341442
rect 135214 341430 135392 341436
rect 130870 341420 131172 341426
rect 130870 341414 131120 341420
rect 135226 341414 135392 341430
rect 135456 341426 135484 341498
rect 135548 341426 135576 341566
rect 137218 341426 137600 341442
rect 139334 341426 139624 341442
rect 139964 341426 139992 341566
rect 164146 341527 164202 341536
rect 164160 341426 164188 341527
rect 164804 341426 164832 341770
rect 316040 341488 316092 341494
rect 288544 341426 288834 341442
rect 290568 341426 290950 341442
rect 292776 341426 293066 341442
rect 296916 341426 297206 341442
rect 299032 341426 299322 341442
rect 322202 341456 322258 341465
rect 316092 341436 316158 341442
rect 316040 341430 316158 341436
rect 135444 341420 135496 341426
rect 131120 341362 131172 341368
rect 135444 341362 135496 341368
rect 135536 341420 135588 341426
rect 137218 341420 137612 341426
rect 137218 341414 137560 341420
rect 135536 341362 135588 341368
rect 139334 341420 139636 341426
rect 139334 341414 139584 341420
rect 137560 341362 137612 341368
rect 139584 341362 139636 341368
rect 139952 341420 140004 341426
rect 139952 341362 140004 341368
rect 164148 341420 164200 341426
rect 164148 341362 164200 341368
rect 164792 341420 164844 341426
rect 164792 341362 164844 341368
rect 288532 341420 288834 341426
rect 288584 341414 288834 341420
rect 290556 341420 290950 341426
rect 288532 341362 288584 341368
rect 290608 341414 290950 341420
rect 292764 341420 293066 341426
rect 290556 341362 290608 341368
rect 292816 341414 293066 341420
rect 296904 341420 297206 341426
rect 292764 341362 292816 341368
rect 296956 341414 297206 341420
rect 299020 341420 299322 341426
rect 296904 341362 296956 341368
rect 299072 341414 299322 341420
rect 316052 341414 316158 341430
rect 326434 341456 326490 341465
rect 322258 341414 322506 341442
rect 322202 341391 322258 341400
rect 328458 341456 328514 341465
rect 326490 341414 326738 341442
rect 326434 341391 326490 341400
rect 330666 341456 330722 341465
rect 328514 341414 328854 341442
rect 328458 341391 328514 341400
rect 330722 341414 330970 341442
rect 330666 341391 330722 341400
rect 299020 341362 299072 341368
rect 331876 272542 331904 344286
rect 331968 272610 331996 344354
rect 577596 343800 577648 343806
rect 577596 343742 577648 343748
rect 577504 343732 577556 343738
rect 577504 343674 577556 343680
rect 331956 272604 332008 272610
rect 331956 272546 332008 272552
rect 331864 272536 331916 272542
rect 331864 272478 331916 272484
rect 92216 97986 92244 102068
rect 92480 99884 92532 99890
rect 92480 99826 92532 99832
rect 92204 97980 92256 97986
rect 92204 97922 92256 97928
rect 92112 20664 92164 20670
rect 92112 20606 92164 20612
rect 91100 7676 91152 7682
rect 91100 7618 91152 7624
rect 91560 7676 91612 7682
rect 91560 7618 91612 7624
rect 87972 7404 88024 7410
rect 87972 7346 88024 7352
rect 86868 4684 86920 4690
rect 86868 4626 86920 4632
rect 86880 480 86908 4626
rect 87984 480 88012 7346
rect 90364 4616 90416 4622
rect 90364 4558 90416 4564
rect 89168 3256 89220 3262
rect 89168 3198 89220 3204
rect 89180 480 89208 3198
rect 90376 480 90404 4558
rect 91572 480 91600 7618
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 78558 -960 78670 326
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92492 354 92520 99826
rect 92676 98002 92704 102037
rect 92572 97980 92624 97986
rect 92676 97974 92796 98002
rect 92572 97922 92624 97928
rect 92584 4826 92612 97922
rect 92664 97912 92716 97918
rect 92664 97854 92716 97860
rect 92676 7750 92704 97854
rect 92664 7744 92716 7750
rect 92664 7686 92716 7692
rect 92768 7614 92796 97974
rect 93136 97918 93164 102037
rect 93596 97986 93624 102037
rect 93860 99748 93912 99754
rect 93860 99690 93912 99696
rect 93584 97980 93636 97986
rect 93584 97922 93636 97928
rect 93124 97912 93176 97918
rect 93124 97854 93176 97860
rect 92756 7608 92808 7614
rect 92756 7550 92808 7556
rect 92572 4820 92624 4826
rect 92572 4762 92624 4768
rect 93872 3466 93900 99690
rect 94148 99634 94176 102037
rect 94608 99754 94636 102037
rect 94596 99748 94648 99754
rect 94596 99690 94648 99696
rect 93964 99606 94176 99634
rect 93964 6914 93992 99606
rect 95068 84194 95096 102037
rect 95620 98002 95648 102037
rect 96080 100026 96108 102037
rect 96068 100020 96120 100026
rect 96068 99962 96120 99968
rect 94056 84166 95096 84194
rect 95344 97974 95648 98002
rect 94056 7818 94084 84166
rect 94044 7812 94096 7818
rect 94044 7754 94096 7760
rect 93964 6886 94084 6914
rect 93952 4820 94004 4826
rect 93952 4762 94004 4768
rect 93860 3460 93912 3466
rect 93860 3402 93912 3408
rect 93964 480 93992 4762
rect 94056 3369 94084 6886
rect 95148 5976 95200 5982
rect 95148 5918 95200 5924
rect 94042 3360 94098 3369
rect 94042 3295 94098 3304
rect 95160 480 95188 5918
rect 95344 4894 95372 97974
rect 96540 84194 96568 102037
rect 97000 98002 97028 102037
rect 95436 84166 96568 84194
rect 96632 97974 97028 98002
rect 95332 4888 95384 4894
rect 95332 4830 95384 4836
rect 95436 3602 95464 84166
rect 96632 4962 96660 97974
rect 97552 84194 97580 102037
rect 98012 98002 98040 102037
rect 98012 97974 98132 98002
rect 98000 97912 98052 97918
rect 98000 97854 98052 97860
rect 96724 84166 97580 84194
rect 96724 6225 96752 84166
rect 96710 6216 96766 6225
rect 96710 6151 96766 6160
rect 96620 4956 96672 4962
rect 96620 4898 96672 4904
rect 97448 4888 97500 4894
rect 97448 4830 97500 4836
rect 95424 3596 95476 3602
rect 95424 3538 95476 3544
rect 96252 3460 96304 3466
rect 96252 3402 96304 3408
rect 96264 480 96292 3402
rect 97460 480 97488 4830
rect 98012 3670 98040 97854
rect 98000 3664 98052 3670
rect 98000 3606 98052 3612
rect 98104 3534 98132 97974
rect 98472 97918 98500 102037
rect 98460 97912 98512 97918
rect 98460 97854 98512 97860
rect 99024 84194 99052 102037
rect 99380 99816 99432 99822
rect 99380 99758 99432 99764
rect 98196 84166 99052 84194
rect 98196 5030 98224 84166
rect 98644 7608 98696 7614
rect 98644 7550 98696 7556
rect 98184 5024 98236 5030
rect 98184 4966 98236 4972
rect 98092 3528 98144 3534
rect 98092 3470 98144 3476
rect 98656 480 98684 7550
rect 99392 6914 99420 99758
rect 99484 7886 99512 102037
rect 99944 100230 99972 102037
rect 99932 100224 99984 100230
rect 99932 100166 99984 100172
rect 100404 100094 100432 102037
rect 100392 100088 100444 100094
rect 100392 100030 100444 100036
rect 100956 98002 100984 102037
rect 100760 97980 100812 97986
rect 100760 97922 100812 97928
rect 100864 97974 100984 98002
rect 99472 7880 99524 7886
rect 99472 7822 99524 7828
rect 99392 6886 99880 6914
rect 99852 480 99880 6886
rect 100772 3738 100800 97922
rect 100864 5098 100892 97974
rect 101416 84194 101444 102037
rect 101876 97986 101904 102037
rect 102428 100162 102456 102037
rect 102416 100156 102468 100162
rect 102416 100098 102468 100104
rect 101864 97980 101916 97986
rect 101864 97922 101916 97928
rect 102232 97980 102284 97986
rect 102232 97922 102284 97928
rect 100956 84166 101444 84194
rect 100956 7954 100984 84166
rect 102244 8974 102272 97922
rect 102888 84194 102916 102037
rect 103348 97986 103376 102037
rect 103900 100298 103928 102037
rect 103888 100292 103940 100298
rect 103888 100234 103940 100240
rect 103336 97980 103388 97986
rect 103336 97922 103388 97928
rect 103612 97980 103664 97986
rect 103612 97922 103664 97928
rect 102336 84166 102916 84194
rect 102232 8968 102284 8974
rect 102232 8910 102284 8916
rect 102336 8022 102364 84166
rect 103624 9042 103652 97922
rect 104360 84194 104388 102037
rect 104820 97986 104848 102037
rect 104900 100020 104952 100026
rect 104900 99962 104952 99968
rect 104808 97980 104860 97986
rect 104808 97922 104860 97928
rect 103716 84166 104388 84194
rect 103612 9036 103664 9042
rect 103612 8978 103664 8984
rect 103716 8090 103744 84166
rect 103704 8084 103756 8090
rect 103704 8026 103756 8032
rect 102324 8016 102376 8022
rect 102324 7958 102376 7964
rect 100944 7948 100996 7954
rect 100944 7890 100996 7896
rect 100852 5092 100904 5098
rect 100852 5034 100904 5040
rect 104532 5024 104584 5030
rect 104532 4966 104584 4972
rect 101036 4956 101088 4962
rect 101036 4898 101088 4904
rect 100760 3732 100812 3738
rect 100760 3674 100812 3680
rect 101048 480 101076 4898
rect 102232 3596 102284 3602
rect 102232 3538 102284 3544
rect 102244 480 102272 3538
rect 103336 3528 103388 3534
rect 103336 3470 103388 3476
rect 103348 480 103376 3470
rect 104544 480 104572 4966
rect 104912 3482 104940 99962
rect 105280 97968 105308 102037
rect 105004 97940 105308 97968
rect 105004 3806 105032 97940
rect 105832 84194 105860 102037
rect 106292 97968 106320 102037
rect 106752 100366 106780 102037
rect 106740 100360 106792 100366
rect 106740 100302 106792 100308
rect 106556 100156 106608 100162
rect 106556 100098 106608 100104
rect 106292 97940 106504 97968
rect 106372 97844 106424 97850
rect 106372 97786 106424 97792
rect 106280 97028 106332 97034
rect 106280 96970 106332 96976
rect 105096 84166 105860 84194
rect 105096 8158 105124 84166
rect 105084 8152 105136 8158
rect 105084 8094 105136 8100
rect 104992 3800 105044 3806
rect 104992 3742 105044 3748
rect 104912 3454 105768 3482
rect 105740 480 105768 3454
rect 106292 490 106320 96970
rect 106384 6186 106412 97786
rect 106476 9110 106504 97940
rect 106568 97034 106596 100098
rect 107304 97850 107332 102037
rect 107660 97980 107712 97986
rect 107764 97968 107792 102037
rect 108224 97986 108252 102037
rect 108304 100292 108356 100298
rect 108304 100234 108356 100240
rect 108212 97980 108264 97986
rect 107764 97940 107884 97968
rect 107660 97922 107712 97928
rect 107292 97844 107344 97850
rect 107292 97786 107344 97792
rect 106556 97028 106608 97034
rect 106556 96970 106608 96976
rect 106464 9104 106516 9110
rect 106464 9046 106516 9052
rect 106372 6180 106424 6186
rect 106372 6122 106424 6128
rect 107672 3874 107700 97922
rect 107752 97844 107804 97850
rect 107752 97786 107804 97792
rect 107764 6254 107792 97786
rect 107856 9178 107884 97940
rect 108212 97922 108264 97928
rect 107844 9172 107896 9178
rect 107844 9114 107896 9120
rect 107752 6248 107804 6254
rect 107752 6190 107804 6196
rect 107660 3868 107712 3874
rect 107660 3810 107712 3816
rect 108316 3602 108344 100234
rect 108684 97850 108712 102037
rect 109236 97968 109264 102037
rect 109696 100434 109724 102037
rect 109684 100428 109736 100434
rect 109684 100370 109736 100376
rect 109144 97940 109264 97968
rect 108672 97844 108724 97850
rect 108672 97786 108724 97792
rect 109144 9246 109172 97940
rect 110156 84194 110184 102037
rect 110420 100088 110472 100094
rect 110420 100030 110472 100036
rect 109236 84166 110184 84194
rect 109132 9240 109184 9246
rect 109132 9182 109184 9188
rect 109236 6322 109264 84166
rect 110432 11778 110460 100030
rect 110604 98048 110656 98054
rect 110604 97990 110656 97996
rect 110512 97980 110564 97986
rect 110512 97922 110564 97928
rect 110524 11914 110552 97922
rect 110616 12186 110644 97990
rect 110708 16574 110736 102037
rect 111168 97986 111196 102037
rect 111628 98054 111656 102037
rect 111800 100224 111852 100230
rect 111800 100166 111852 100172
rect 111616 98048 111668 98054
rect 111616 97990 111668 97996
rect 111156 97980 111208 97986
rect 111156 97922 111208 97928
rect 110708 16546 110920 16574
rect 110616 12158 110828 12186
rect 110524 11886 110644 11914
rect 110432 11750 110552 11778
rect 110420 11688 110472 11694
rect 110420 11630 110472 11636
rect 109224 6316 109276 6322
rect 109224 6258 109276 6264
rect 110432 3942 110460 11630
rect 110420 3936 110472 3942
rect 110420 3878 110472 3884
rect 108304 3596 108356 3602
rect 108304 3538 108356 3544
rect 109314 3360 109370 3369
rect 109314 3295 109370 3304
rect 108120 2848 108172 2854
rect 108120 2790 108172 2796
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106292 462 106504 490
rect 108132 480 108160 2790
rect 109328 480 109356 3295
rect 110524 480 110552 11750
rect 110616 11694 110644 11886
rect 110604 11688 110656 11694
rect 110604 11630 110656 11636
rect 110800 8226 110828 12158
rect 110892 9314 110920 16546
rect 110880 9308 110932 9314
rect 110880 9250 110932 9256
rect 110788 8220 110840 8226
rect 110788 8162 110840 8168
rect 111616 3732 111668 3738
rect 111616 3674 111668 3680
rect 111628 480 111656 3674
rect 111812 490 111840 100166
rect 112088 97968 112116 102037
rect 112640 100502 112668 102037
rect 112628 100496 112680 100502
rect 112628 100438 112680 100444
rect 111904 97940 112116 97968
rect 111904 6390 111932 97940
rect 113100 84194 113128 102037
rect 113180 97980 113232 97986
rect 113180 97922 113232 97928
rect 111996 84166 113128 84194
rect 111996 8294 112024 84166
rect 111984 8288 112036 8294
rect 111984 8230 112036 8236
rect 111892 6384 111944 6390
rect 111892 6326 111944 6332
rect 113192 4010 113220 97922
rect 113560 84194 113588 102037
rect 114112 97986 114140 102037
rect 114100 97980 114152 97986
rect 114100 97922 114152 97928
rect 114572 93854 114600 102037
rect 114572 93826 114692 93854
rect 113284 84166 113588 84194
rect 113284 6458 113312 84166
rect 114664 7546 114692 93826
rect 115032 84194 115060 102037
rect 115584 100570 115612 102037
rect 115572 100564 115624 100570
rect 115572 100506 115624 100512
rect 115940 100360 115992 100366
rect 115940 100302 115992 100308
rect 114756 84166 115060 84194
rect 114652 7540 114704 7546
rect 114652 7482 114704 7488
rect 114756 6526 114784 84166
rect 114744 6520 114796 6526
rect 114744 6462 114796 6468
rect 113272 6452 113324 6458
rect 113272 6394 113324 6400
rect 115204 4548 115256 4554
rect 115204 4490 115256 4496
rect 113180 4004 113232 4010
rect 113180 3946 113232 3952
rect 114008 3596 114060 3602
rect 114008 3538 114060 3544
rect 106476 354 106504 462
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 111812 462 112392 490
rect 114020 480 114048 3538
rect 115216 2854 115244 4490
rect 115952 3482 115980 100302
rect 116044 98002 116072 102037
rect 116044 97974 116164 98002
rect 116032 97912 116084 97918
rect 116032 97854 116084 97860
rect 116044 4078 116072 97854
rect 116136 5166 116164 97974
rect 116504 84194 116532 102037
rect 116964 97918 116992 102037
rect 117320 100496 117372 100502
rect 117320 100438 117372 100444
rect 116952 97912 117004 97918
rect 116952 97854 117004 97860
rect 116228 84166 116532 84194
rect 116228 6594 116256 84166
rect 116216 6588 116268 6594
rect 116216 6530 116268 6536
rect 116124 5160 116176 5166
rect 116124 5102 116176 5108
rect 117228 5160 117280 5166
rect 117228 5102 117280 5108
rect 116032 4072 116084 4078
rect 116032 4014 116084 4020
rect 117240 3738 117268 5102
rect 117228 3732 117280 3738
rect 117228 3674 117280 3680
rect 115952 3454 116440 3482
rect 115204 2848 115256 2854
rect 115204 2790 115256 2796
rect 115296 2848 115348 2854
rect 115296 2790 115348 2796
rect 115308 2530 115336 2790
rect 115216 2502 115336 2530
rect 115216 480 115244 2502
rect 116412 480 116440 3454
rect 112364 354 112392 462
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117332 354 117360 100438
rect 117516 98002 117544 102037
rect 117424 97974 117544 98002
rect 117424 5234 117452 97974
rect 117976 84194 118004 102037
rect 118436 100638 118464 102037
rect 118424 100632 118476 100638
rect 118424 100574 118476 100580
rect 118988 98002 119016 102037
rect 118700 97980 118752 97986
rect 118700 97922 118752 97928
rect 118804 97974 119016 98002
rect 117516 84166 118004 84194
rect 117516 6662 117544 84166
rect 117504 6656 117556 6662
rect 117504 6598 117556 6604
rect 117412 5228 117464 5234
rect 117412 5170 117464 5176
rect 118608 5092 118660 5098
rect 118608 5034 118660 5040
rect 118620 2854 118648 5034
rect 118712 4146 118740 97922
rect 118804 4865 118832 97974
rect 119448 84194 119476 102037
rect 119908 97986 119936 102037
rect 119896 97980 119948 97986
rect 119896 97922 119948 97928
rect 120172 97980 120224 97986
rect 120172 97922 120224 97928
rect 118896 84166 119476 84194
rect 118896 6730 118924 84166
rect 120184 6798 120212 97922
rect 120368 84194 120396 102037
rect 120920 97986 120948 102037
rect 121380 100706 121408 102037
rect 121368 100700 121420 100706
rect 121368 100642 121420 100648
rect 121460 100428 121512 100434
rect 121460 100370 121512 100376
rect 120908 97980 120960 97986
rect 120908 97922 120960 97928
rect 120276 84166 120396 84194
rect 120172 6792 120224 6798
rect 120172 6734 120224 6740
rect 118884 6724 118936 6730
rect 118884 6666 118936 6672
rect 120276 5302 120304 84166
rect 120264 5296 120316 5302
rect 120264 5238 120316 5244
rect 118790 4856 118846 4865
rect 118790 4791 118846 4800
rect 118700 4140 118752 4146
rect 118700 4082 118752 4088
rect 121092 3800 121144 3806
rect 121092 3742 121144 3748
rect 119896 3732 119948 3738
rect 119896 3674 119948 3680
rect 118792 3664 118844 3670
rect 118792 3606 118844 3612
rect 118608 2848 118660 2854
rect 118608 2790 118660 2796
rect 118804 480 118832 3606
rect 119908 480 119936 3674
rect 121104 480 121132 3742
rect 121472 3482 121500 100370
rect 121840 98002 121868 102037
rect 121564 97974 121868 98002
rect 121564 5370 121592 97974
rect 122392 84194 122420 102037
rect 121656 84166 122420 84194
rect 121656 6866 121684 84166
rect 121644 6860 121696 6866
rect 121644 6802 121696 6808
rect 121552 5364 121604 5370
rect 121552 5306 121604 5312
rect 121472 3454 122328 3482
rect 122300 480 122328 3454
rect 122852 3398 122880 102037
rect 123312 98002 123340 102037
rect 122944 97974 123340 98002
rect 122944 5438 122972 97974
rect 123772 84194 123800 102037
rect 124324 99958 124352 102037
rect 124312 99952 124364 99958
rect 124312 99894 124364 99900
rect 124784 98138 124812 102037
rect 123036 84166 123800 84194
rect 124324 98110 124812 98138
rect 123036 6118 123064 84166
rect 123024 6112 123076 6118
rect 123024 6054 123076 6060
rect 124324 5506 124352 98110
rect 125244 98002 125272 102037
rect 125324 100564 125376 100570
rect 125324 100506 125376 100512
rect 124416 97974 125272 98002
rect 124416 6050 124444 97974
rect 125336 84194 125364 100506
rect 125796 98002 125824 102037
rect 124508 84166 125364 84194
rect 125612 97974 125824 98002
rect 124508 16574 124536 84166
rect 124508 16546 124720 16574
rect 124404 6044 124456 6050
rect 124404 5986 124456 5992
rect 124312 5500 124364 5506
rect 124312 5442 124364 5448
rect 122932 5432 122984 5438
rect 122932 5374 122984 5380
rect 123484 3868 123536 3874
rect 123484 3810 123536 3816
rect 122840 3392 122892 3398
rect 122840 3334 122892 3340
rect 123496 480 123524 3810
rect 124692 480 124720 16546
rect 125612 3330 125640 97974
rect 126256 97866 126284 102037
rect 125704 97838 126284 97866
rect 125704 4758 125732 97838
rect 126716 84194 126744 102037
rect 127072 98048 127124 98054
rect 127072 97990 127124 97996
rect 126980 97980 127032 97986
rect 126980 97922 127032 97928
rect 125796 84166 126744 84194
rect 125796 7478 125824 84166
rect 125784 7472 125836 7478
rect 125784 7414 125836 7420
rect 125692 4752 125744 4758
rect 125692 4694 125744 4700
rect 126992 4690 127020 97922
rect 127084 7410 127112 97990
rect 127268 84194 127296 102037
rect 127728 97986 127756 102037
rect 128188 98054 128216 102037
rect 128176 98048 128228 98054
rect 128648 98002 128676 102037
rect 128176 97990 128228 97996
rect 127716 97980 127768 97986
rect 127716 97922 127768 97928
rect 128372 97974 128676 98002
rect 127176 84166 127296 84194
rect 127176 9382 127204 84166
rect 127164 9376 127216 9382
rect 127164 9318 127216 9324
rect 127072 7404 127124 7410
rect 127072 7346 127124 7352
rect 126980 4684 127032 4690
rect 126980 4626 127032 4632
rect 126980 4004 127032 4010
rect 126980 3946 127032 3952
rect 125876 3936 125928 3942
rect 125876 3878 125928 3884
rect 125600 3324 125652 3330
rect 125600 3266 125652 3272
rect 125888 480 125916 3878
rect 126992 480 127020 3946
rect 128372 3262 128400 97974
rect 129200 97866 129228 102037
rect 129280 100632 129332 100638
rect 129280 100574 129332 100580
rect 128464 97838 129228 97866
rect 128464 4622 128492 97838
rect 128544 97776 128596 97782
rect 128544 97718 128596 97724
rect 128556 7682 128584 97718
rect 129292 84194 129320 100574
rect 129660 97782 129688 102037
rect 130120 99890 130148 102037
rect 130108 99884 130160 99890
rect 130108 99826 130160 99832
rect 129648 97776 129700 97782
rect 129648 97718 129700 97724
rect 130672 84194 130700 102037
rect 131132 99770 131160 102037
rect 131132 99742 131344 99770
rect 131120 98048 131172 98054
rect 131120 97990 131172 97996
rect 129016 84166 129320 84194
rect 129844 84166 130700 84194
rect 128544 7676 128596 7682
rect 128544 7618 128596 7624
rect 128452 4616 128504 4622
rect 128452 4558 128504 4564
rect 128360 3256 128412 3262
rect 128360 3198 128412 3204
rect 129016 3058 129044 84166
rect 129844 4826 129872 84166
rect 129832 4820 129884 4826
rect 129832 4762 129884 4768
rect 130568 4140 130620 4146
rect 130568 4082 130620 4088
rect 129372 4072 129424 4078
rect 129372 4014 129424 4020
rect 128176 3052 128228 3058
rect 128176 2994 128228 3000
rect 129004 3052 129056 3058
rect 129004 2994 129056 3000
rect 128188 480 128216 2994
rect 129384 480 129412 4014
rect 130580 480 130608 4082
rect 131132 3466 131160 97990
rect 131212 97980 131264 97986
rect 131212 97922 131264 97928
rect 131224 4894 131252 97922
rect 131316 5982 131344 99742
rect 131592 98054 131620 102037
rect 131580 98048 131632 98054
rect 131580 97990 131632 97996
rect 132052 97986 132080 102037
rect 132040 97980 132092 97986
rect 132040 97922 132092 97928
rect 132604 7614 132632 102037
rect 133064 99822 133092 102037
rect 133052 99816 133104 99822
rect 133052 99758 133104 99764
rect 133524 84194 133552 102037
rect 134076 100298 134104 102037
rect 134064 100292 134116 100298
rect 134064 100234 134116 100240
rect 133972 98184 134024 98190
rect 133972 98126 134024 98132
rect 132696 84166 133552 84194
rect 132592 7608 132644 7614
rect 132592 7550 132644 7556
rect 131304 5976 131356 5982
rect 131304 5918 131356 5924
rect 132696 4962 132724 84166
rect 133984 5030 134012 98126
rect 134536 84194 134564 102037
rect 134996 98190 135024 102037
rect 135456 100026 135484 102037
rect 136008 100162 136036 102037
rect 135996 100156 136048 100162
rect 135996 100098 136048 100104
rect 135444 100020 135496 100026
rect 135444 99962 135496 99968
rect 134984 98184 135036 98190
rect 134984 98126 135036 98132
rect 136468 84194 136496 102037
rect 136928 98002 136956 102037
rect 137008 100292 137060 100298
rect 137008 100234 137060 100240
rect 134076 84166 134564 84194
rect 135364 84166 136496 84194
rect 136744 97974 136956 98002
rect 133972 5024 134024 5030
rect 133972 4966 134024 4972
rect 132684 4956 132736 4962
rect 132684 4898 132736 4904
rect 131212 4888 131264 4894
rect 131212 4830 131264 4836
rect 134076 3534 134104 84166
rect 135364 4554 135392 84166
rect 135352 4548 135404 4554
rect 135352 4490 135404 4496
rect 134064 3528 134116 3534
rect 134064 3470 134116 3476
rect 135260 3528 135312 3534
rect 135260 3470 135312 3476
rect 131120 3460 131172 3466
rect 131120 3402 131172 3408
rect 132960 3460 133012 3466
rect 132960 3402 133012 3408
rect 131764 3392 131816 3398
rect 131764 3334 131816 3340
rect 131776 480 131804 3334
rect 132972 480 133000 3402
rect 134156 3256 134208 3262
rect 134156 3198 134208 3204
rect 134168 480 134196 3198
rect 135272 480 135300 3470
rect 136744 3369 136772 97974
rect 136824 97912 136876 97918
rect 136824 97854 136876 97860
rect 136836 5166 136864 97854
rect 137020 84194 137048 100234
rect 137480 100094 137508 102037
rect 137468 100088 137520 100094
rect 137468 100030 137520 100036
rect 137940 97918 137968 102037
rect 138400 100230 138428 102037
rect 138388 100224 138440 100230
rect 138388 100166 138440 100172
rect 138020 100020 138072 100026
rect 138020 99962 138072 99968
rect 137928 97912 137980 97918
rect 137928 97854 137980 97860
rect 136928 84166 137048 84194
rect 136928 16574 136956 84166
rect 136928 16546 137232 16574
rect 136824 5160 136876 5166
rect 136824 5102 136876 5108
rect 136730 3360 136786 3369
rect 136456 3324 136508 3330
rect 136730 3295 136786 3304
rect 136456 3266 136508 3272
rect 136468 480 136496 3266
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 138032 3482 138060 99962
rect 138952 84194 138980 102037
rect 139412 100314 139440 102037
rect 139872 100366 139900 102037
rect 140332 100502 140360 102037
rect 140320 100496 140372 100502
rect 140320 100438 140372 100444
rect 139860 100360 139912 100366
rect 139412 100286 139716 100314
rect 139860 100302 139912 100308
rect 139400 100156 139452 100162
rect 139400 100098 139452 100104
rect 138124 84166 138980 84194
rect 138124 3602 138152 84166
rect 138112 3596 138164 3602
rect 138112 3538 138164 3544
rect 138032 3454 138888 3482
rect 138860 480 138888 3454
rect 139412 490 139440 100098
rect 139688 96914 139716 100286
rect 140884 98002 140912 102037
rect 140780 97980 140832 97986
rect 140884 97974 141004 98002
rect 140780 97922 140832 97928
rect 139504 96886 139716 96914
rect 139504 5098 139532 96886
rect 139492 5092 139544 5098
rect 139492 5034 139544 5040
rect 140792 3806 140820 97922
rect 140872 97912 140924 97918
rect 140872 97854 140924 97860
rect 140780 3800 140832 3806
rect 140780 3742 140832 3748
rect 140884 3738 140912 97854
rect 140872 3732 140924 3738
rect 140872 3674 140924 3680
rect 140976 3670 141004 97974
rect 141344 97918 141372 102037
rect 141804 97986 141832 102037
rect 142356 100434 142384 102037
rect 142344 100428 142396 100434
rect 142344 100370 142396 100376
rect 141792 97980 141844 97986
rect 141792 97922 141844 97928
rect 141332 97912 141384 97918
rect 141332 97854 141384 97860
rect 142816 84194 142844 102037
rect 143276 100570 143304 102037
rect 143264 100564 143316 100570
rect 143264 100506 143316 100512
rect 143540 99612 143592 99618
rect 143540 99554 143592 99560
rect 142264 84166 142844 84194
rect 142264 3874 142292 84166
rect 142252 3868 142304 3874
rect 142252 3810 142304 3816
rect 142436 3800 142488 3806
rect 142436 3742 142488 3748
rect 140964 3664 141016 3670
rect 140964 3606 141016 3612
rect 141240 3664 141292 3670
rect 141240 3606 141292 3612
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139412 462 139624 490
rect 141252 480 141280 3606
rect 142448 480 142476 3742
rect 143552 480 143580 99554
rect 143632 97980 143684 97986
rect 143632 97922 143684 97928
rect 143644 4010 143672 97922
rect 143632 4004 143684 4010
rect 143632 3946 143684 3952
rect 143736 3942 143764 102037
rect 144288 97986 144316 102037
rect 144748 100638 144776 102037
rect 144736 100632 144788 100638
rect 144736 100574 144788 100580
rect 144276 97980 144328 97986
rect 144276 97922 144328 97928
rect 144920 97980 144972 97986
rect 145208 97968 145236 102037
rect 145760 97986 145788 102037
rect 144920 97922 144972 97928
rect 145024 97940 145236 97968
rect 145748 97980 145800 97986
rect 144932 4146 144960 97922
rect 144920 4140 144972 4146
rect 144920 4082 144972 4088
rect 145024 4078 145052 97940
rect 145748 97922 145800 97928
rect 146220 84194 146248 102037
rect 146300 100632 146352 100638
rect 146300 100574 146352 100580
rect 145116 84166 146248 84194
rect 145012 4072 145064 4078
rect 145012 4014 145064 4020
rect 143724 3936 143776 3942
rect 143724 3878 143776 3884
rect 145116 3398 145144 84166
rect 145104 3392 145156 3398
rect 145104 3334 145156 3340
rect 145932 3120 145984 3126
rect 146312 3108 146340 100574
rect 146392 97980 146444 97986
rect 146392 97922 146444 97928
rect 146404 3262 146432 97922
rect 146680 84194 146708 102037
rect 147232 97986 147260 102037
rect 147692 99374 147720 102037
rect 147692 99346 147904 99374
rect 147220 97980 147272 97986
rect 147220 97922 147272 97928
rect 147772 94580 147824 94586
rect 147772 94522 147824 94528
rect 146496 84166 146708 84194
rect 146496 3602 146524 84166
rect 146484 3596 146536 3602
rect 146484 3538 146536 3544
rect 147784 3330 147812 94522
rect 147876 3670 147904 99346
rect 148152 94586 148180 102037
rect 148612 100298 148640 102037
rect 148600 100292 148652 100298
rect 148600 100234 148652 100240
rect 148232 100224 148284 100230
rect 148232 100166 148284 100172
rect 148140 94580 148192 94586
rect 148140 94522 148192 94528
rect 148244 84194 148272 100166
rect 149164 100026 149192 102037
rect 149624 100162 149652 102037
rect 149612 100156 149664 100162
rect 149612 100098 149664 100104
rect 149152 100020 149204 100026
rect 149152 99962 149204 99968
rect 150084 84194 150112 102037
rect 150532 94580 150584 94586
rect 150532 94522 150584 94528
rect 147968 84166 148272 84194
rect 149164 84166 150112 84194
rect 147864 3664 147916 3670
rect 147864 3606 147916 3612
rect 147772 3324 147824 3330
rect 147772 3266 147824 3272
rect 146392 3256 146444 3262
rect 146392 3198 146444 3204
rect 146312 3080 147168 3108
rect 145932 3062 145984 3068
rect 144736 3052 144788 3058
rect 144736 2994 144788 3000
rect 144748 480 144776 2994
rect 145944 480 145972 3062
rect 147140 480 147168 3080
rect 139596 354 139624 462
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 147968 354 147996 84166
rect 149164 3738 149192 84166
rect 149152 3732 149204 3738
rect 149152 3674 149204 3680
rect 150544 3058 150572 94522
rect 150636 3806 150664 102037
rect 150716 100020 150768 100026
rect 150716 99962 150768 99968
rect 150624 3800 150676 3806
rect 150624 3742 150676 3748
rect 150728 3482 150756 99962
rect 151096 99618 151124 102037
rect 151084 99612 151136 99618
rect 151084 99554 151136 99560
rect 151556 94586 151584 102037
rect 151820 100292 151872 100298
rect 151820 100234 151872 100240
rect 151544 94580 151596 94586
rect 151544 94522 151596 94528
rect 150636 3454 150756 3482
rect 150532 3052 150584 3058
rect 150532 2994 150584 3000
rect 149520 2984 149572 2990
rect 149520 2926 149572 2932
rect 149532 480 149560 2926
rect 150636 480 150664 3454
rect 151832 480 151860 100234
rect 152016 84194 152044 102037
rect 152568 100638 152596 102037
rect 152556 100632 152608 100638
rect 152556 100574 152608 100580
rect 153028 100230 153056 102037
rect 153016 100224 153068 100230
rect 153016 100166 153068 100172
rect 153488 84194 153516 102037
rect 154040 100026 154068 102037
rect 154500 100298 154528 102037
rect 154488 100292 154540 100298
rect 154488 100234 154540 100240
rect 154028 100020 154080 100026
rect 154028 99962 154080 99968
rect 154580 94580 154632 94586
rect 154580 94522 154632 94528
rect 151924 84166 152044 84194
rect 153396 84166 153516 84194
rect 151924 3126 151952 84166
rect 153016 3528 153068 3534
rect 153016 3470 153068 3476
rect 151912 3120 151964 3126
rect 151912 3062 151964 3068
rect 153028 480 153056 3470
rect 153396 2990 153424 84166
rect 154592 3482 154620 94522
rect 154960 84194 154988 102037
rect 155420 94586 155448 102037
rect 155972 99374 156000 102037
rect 155972 99346 156092 99374
rect 155408 94580 155460 94586
rect 155408 94522 155460 94528
rect 155960 94580 156012 94586
rect 155960 94522 156012 94528
rect 154684 84166 154988 84194
rect 154684 3534 154712 84166
rect 155972 3534 156000 94522
rect 154224 3454 154620 3482
rect 154672 3528 154724 3534
rect 154672 3470 154724 3476
rect 155960 3528 156012 3534
rect 155960 3470 156012 3476
rect 153384 2984 153436 2990
rect 153384 2926 153436 2932
rect 154224 480 154252 3454
rect 156064 2802 156092 99346
rect 156432 94586 156460 102037
rect 156892 100502 156920 102037
rect 157444 100570 157472 102037
rect 157432 100564 157484 100570
rect 157432 100506 157484 100512
rect 156880 100496 156932 100502
rect 156880 100438 156932 100444
rect 157340 100496 157392 100502
rect 157340 100438 157392 100444
rect 156420 94580 156472 94586
rect 156420 94522 156472 94528
rect 156236 3528 156288 3534
rect 156236 3470 156288 3476
rect 157352 3482 157380 100438
rect 157904 98002 157932 102037
rect 157444 97974 157932 98002
rect 157444 3670 157472 97974
rect 158364 84194 158392 102037
rect 158720 100564 158772 100570
rect 158720 100506 158772 100512
rect 157536 84166 158392 84194
rect 157536 3738 157564 84166
rect 157524 3732 157576 3738
rect 157524 3674 157576 3680
rect 157432 3664 157484 3670
rect 157432 3606 157484 3612
rect 158732 3482 158760 100506
rect 158916 100366 158944 102037
rect 158904 100360 158956 100366
rect 158904 100302 158956 100308
rect 158812 98524 158864 98530
rect 158812 98466 158864 98472
rect 158824 3602 158852 98466
rect 159376 84194 159404 102037
rect 159836 98530 159864 102037
rect 160296 100026 160324 102037
rect 160284 100020 160336 100026
rect 160284 99962 160336 99968
rect 159824 98524 159876 98530
rect 159824 98466 159876 98472
rect 160100 97980 160152 97986
rect 160100 97922 160152 97928
rect 158916 84166 159404 84194
rect 158916 16574 158944 84166
rect 158916 16546 159036 16574
rect 159008 4146 159036 16546
rect 158996 4140 159048 4146
rect 158996 4082 159048 4088
rect 160112 4078 160140 97922
rect 160848 84194 160876 102037
rect 161308 97986 161336 102037
rect 161572 101856 161624 101862
rect 161572 101798 161624 101804
rect 161480 100360 161532 100366
rect 161480 100302 161532 100308
rect 161296 97980 161348 97986
rect 161296 97922 161348 97928
rect 160204 84166 160876 84194
rect 160100 4072 160152 4078
rect 160100 4014 160152 4020
rect 160100 3664 160152 3670
rect 160100 3606 160152 3612
rect 158812 3596 158864 3602
rect 158812 3538 158864 3544
rect 155880 2774 156092 2802
rect 148294 354 148406 480
rect 147968 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 354 155490 480
rect 155880 354 155908 2774
rect 155378 326 155908 354
rect 156248 354 156276 3470
rect 157352 3454 157840 3482
rect 158732 3454 158944 3482
rect 157812 480 157840 3454
rect 158916 480 158944 3454
rect 160112 480 160140 3606
rect 160204 3466 160232 84166
rect 161296 3732 161348 3738
rect 161296 3674 161348 3680
rect 160192 3460 160244 3466
rect 160192 3402 160244 3408
rect 161308 480 161336 3674
rect 161492 490 161520 100302
rect 161584 4010 161612 101798
rect 161768 84194 161796 102037
rect 162320 99550 162348 102037
rect 162780 101862 162808 102037
rect 162768 101856 162820 101862
rect 162768 101798 162820 101804
rect 162308 99544 162360 99550
rect 162308 99486 162360 99492
rect 163240 97968 163268 102037
rect 161676 84166 161796 84194
rect 162872 97940 163268 97968
rect 161572 4004 161624 4010
rect 161572 3946 161624 3952
rect 161676 3398 161704 84166
rect 162872 3942 162900 97940
rect 163700 84194 163728 102037
rect 164252 100162 164280 102037
rect 164240 100156 164292 100162
rect 164240 100098 164292 100104
rect 164712 84194 164740 102037
rect 165172 100094 165200 102037
rect 165160 100088 165212 100094
rect 165160 100030 165212 100036
rect 165724 100026 165752 102037
rect 164884 100020 164936 100026
rect 164884 99962 164936 99968
rect 165712 100020 165764 100026
rect 165712 99962 165764 99968
rect 162964 84166 163728 84194
rect 164252 84166 164740 84194
rect 162860 3936 162912 3942
rect 162860 3878 162912 3884
rect 162964 3874 162992 84166
rect 163688 4140 163740 4146
rect 163688 4082 163740 4088
rect 162952 3868 163004 3874
rect 162952 3810 163004 3816
rect 161664 3392 161716 3398
rect 161664 3334 161716 3340
rect 156574 354 156686 480
rect 156248 326 156686 354
rect 155378 -960 155490 326
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 161492 462 162072 490
rect 163700 480 163728 4082
rect 164252 3806 164280 84166
rect 164240 3800 164292 3806
rect 164240 3742 164292 3748
rect 164896 3534 164924 99962
rect 165620 99952 165672 99958
rect 165620 99894 165672 99900
rect 165632 3670 165660 99894
rect 166184 84194 166212 102037
rect 166644 99958 166672 102037
rect 167104 100366 167132 102037
rect 167092 100360 167144 100366
rect 167092 100302 167144 100308
rect 167656 100230 167684 102037
rect 167644 100224 167696 100230
rect 167644 100166 167696 100172
rect 166632 99952 166684 99958
rect 166632 99894 166684 99900
rect 168116 84194 168144 102037
rect 168576 99890 168604 102037
rect 168564 99884 168616 99890
rect 168564 99826 168616 99832
rect 168380 99272 168432 99278
rect 168380 99214 168432 99220
rect 165724 84166 166212 84194
rect 167012 84166 168144 84194
rect 165724 3738 165752 84166
rect 165712 3732 165764 3738
rect 165712 3674 165764 3680
rect 165620 3664 165672 3670
rect 165620 3606 165672 3612
rect 167012 3602 167040 84166
rect 168392 5250 168420 99214
rect 169128 84194 169156 102037
rect 169588 99278 169616 102037
rect 170048 100434 170076 102037
rect 170036 100428 170088 100434
rect 170036 100370 170088 100376
rect 169760 99544 169812 99550
rect 169760 99486 169812 99492
rect 169576 99272 169628 99278
rect 169576 99214 169628 99220
rect 168484 84166 169156 84194
rect 168484 5438 168512 84166
rect 168472 5432 168524 5438
rect 168472 5374 168524 5380
rect 168392 5222 168512 5250
rect 168380 4072 168432 4078
rect 168380 4014 168432 4020
rect 167000 3596 167052 3602
rect 167000 3538 167052 3544
rect 164516 3528 164568 3534
rect 164516 3470 164568 3476
rect 164884 3528 164936 3534
rect 164884 3470 164936 3476
rect 166080 3528 166132 3534
rect 166080 3470 166132 3476
rect 162044 354 162072 462
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164528 354 164556 3470
rect 166092 480 166120 3470
rect 167184 3460 167236 3466
rect 167184 3402 167236 3408
rect 167196 480 167224 3402
rect 168392 480 168420 4014
rect 168484 3534 168512 5222
rect 168472 3528 168524 3534
rect 168472 3470 168524 3476
rect 169576 3392 169628 3398
rect 169576 3334 169628 3340
rect 169588 480 169616 3334
rect 169772 490 169800 99486
rect 169852 97980 169904 97986
rect 169852 97922 169904 97928
rect 169864 3466 169892 97922
rect 170600 84194 170628 102037
rect 171060 97986 171088 102037
rect 171520 100706 171548 102037
rect 171508 100700 171560 100706
rect 171508 100642 171560 100648
rect 171048 97980 171100 97986
rect 171048 97922 171100 97928
rect 171980 84194 172008 102037
rect 169956 84166 170628 84194
rect 171152 84166 172008 84194
rect 169956 5370 169984 84166
rect 169944 5364 169996 5370
rect 169944 5306 169996 5312
rect 171152 5302 171180 84166
rect 171140 5296 171192 5302
rect 171140 5238 171192 5244
rect 172532 4146 172560 102037
rect 172992 100570 173020 102037
rect 172980 100564 173032 100570
rect 172980 100506 173032 100512
rect 173452 84194 173480 102037
rect 174004 98002 174032 102037
rect 174464 100502 174492 102037
rect 174452 100496 174504 100502
rect 174452 100438 174504 100444
rect 172624 84166 173480 84194
rect 173912 97974 174032 98002
rect 172624 5234 172652 84166
rect 172612 5228 172664 5234
rect 172612 5170 172664 5176
rect 172520 4140 172572 4146
rect 172520 4082 172572 4088
rect 173912 4078 173940 97974
rect 174924 84194 174952 102037
rect 175280 100156 175332 100162
rect 175280 100098 175332 100104
rect 174004 84166 174952 84194
rect 174004 5166 174032 84166
rect 173992 5160 174044 5166
rect 173992 5102 174044 5108
rect 173900 4072 173952 4078
rect 173900 4014 173952 4020
rect 171968 4004 172020 4010
rect 171968 3946 172020 3952
rect 169852 3460 169904 3466
rect 169852 3402 169904 3408
rect 164854 354 164966 480
rect 164528 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 169772 462 170352 490
rect 171980 480 172008 3946
rect 173164 3936 173216 3942
rect 173164 3878 173216 3884
rect 173176 480 173204 3878
rect 174268 3868 174320 3874
rect 174268 3810 174320 3816
rect 174280 480 174308 3810
rect 175292 3482 175320 100098
rect 175384 99958 175412 102037
rect 175936 100162 175964 102037
rect 175924 100156 175976 100162
rect 175924 100098 175976 100104
rect 175372 99952 175424 99958
rect 175372 99894 175424 99900
rect 176396 84194 176424 102037
rect 176856 98002 176884 102037
rect 177408 100638 177436 102037
rect 177396 100632 177448 100638
rect 177396 100574 177448 100580
rect 176936 100088 176988 100094
rect 176936 100030 176988 100036
rect 175384 84166 176424 84194
rect 176764 97974 176884 98002
rect 175384 5098 175412 84166
rect 175372 5092 175424 5098
rect 175372 5034 175424 5040
rect 176764 4010 176792 97974
rect 176844 97912 176896 97918
rect 176844 97854 176896 97860
rect 176856 5030 176884 97854
rect 176948 16574 176976 100030
rect 177868 97918 177896 102037
rect 178040 100020 178092 100026
rect 178040 99962 178092 99968
rect 177856 97912 177908 97918
rect 177856 97854 177908 97860
rect 176948 16546 177896 16574
rect 176844 5024 176896 5030
rect 176844 4966 176896 4972
rect 176752 4004 176804 4010
rect 176752 3946 176804 3952
rect 176660 3800 176712 3806
rect 176660 3742 176712 3748
rect 175292 3454 175504 3482
rect 175476 480 175504 3454
rect 176672 480 176700 3742
rect 177868 480 177896 16546
rect 178052 490 178080 99962
rect 178132 97980 178184 97986
rect 178132 97922 178184 97928
rect 178144 4894 178172 97922
rect 178328 84194 178356 102037
rect 178788 100026 178816 102037
rect 178776 100020 178828 100026
rect 178776 99962 178828 99968
rect 179340 97986 179368 102037
rect 179328 97980 179380 97986
rect 179328 97922 179380 97928
rect 179800 84194 179828 102037
rect 180260 100094 180288 102037
rect 180248 100088 180300 100094
rect 180248 100030 180300 100036
rect 180812 97968 180840 102037
rect 180812 97940 180932 97968
rect 180800 97844 180852 97850
rect 180800 97786 180852 97792
rect 178236 84166 178356 84194
rect 179432 84166 179828 84194
rect 178236 4962 178264 84166
rect 178224 4956 178276 4962
rect 178224 4898 178276 4904
rect 178132 4888 178184 4894
rect 178132 4830 178184 4836
rect 179432 3942 179460 84166
rect 180812 4826 180840 97786
rect 180904 6118 180932 97940
rect 181272 97850 181300 102037
rect 181732 100298 181760 102037
rect 182180 100360 182232 100366
rect 182180 100302 182232 100308
rect 181720 100292 181772 100298
rect 181720 100234 181772 100240
rect 181260 97844 181312 97850
rect 181260 97786 181312 97792
rect 180892 6112 180944 6118
rect 180892 6054 180944 6060
rect 180800 4820 180852 4826
rect 180800 4762 180852 4768
rect 179420 3936 179472 3942
rect 179420 3878 179472 3884
rect 180248 3732 180300 3738
rect 180248 3674 180300 3680
rect 170324 354 170352 462
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178052 462 178632 490
rect 180260 480 180288 3674
rect 181444 3664 181496 3670
rect 181444 3606 181496 3612
rect 181456 480 181484 3606
rect 178604 354 178632 462
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182192 354 182220 100302
rect 182284 97968 182312 102037
rect 182284 97940 182404 97968
rect 182272 97844 182324 97850
rect 182272 97786 182324 97792
rect 182284 3874 182312 97786
rect 182376 4554 182404 97940
rect 182744 97850 182772 102037
rect 183204 100366 183232 102037
rect 183192 100360 183244 100366
rect 183192 100302 183244 100308
rect 183560 100224 183612 100230
rect 183560 100166 183612 100172
rect 182732 97844 182784 97850
rect 182732 97786 182784 97792
rect 182364 4548 182416 4554
rect 182364 4490 182416 4496
rect 182272 3868 182324 3874
rect 182272 3810 182324 3816
rect 183572 3482 183600 100166
rect 183664 97968 183692 102037
rect 183664 97940 183784 97968
rect 183652 97844 183704 97850
rect 183652 97786 183704 97792
rect 183664 4622 183692 97786
rect 183756 16574 183784 97940
rect 184216 97850 184244 102037
rect 184676 100230 184704 102037
rect 184664 100224 184716 100230
rect 184664 100166 184716 100172
rect 185032 98116 185084 98122
rect 185032 98058 185084 98064
rect 184204 97844 184256 97850
rect 184204 97786 184256 97792
rect 183756 16546 183876 16574
rect 183848 6186 183876 16546
rect 185044 6866 185072 98058
rect 185032 6860 185084 6866
rect 185032 6802 185084 6808
rect 185136 6798 185164 102037
rect 185308 99884 185360 99890
rect 185308 99826 185360 99832
rect 185216 97980 185268 97986
rect 185216 97922 185268 97928
rect 185124 6792 185176 6798
rect 185124 6734 185176 6740
rect 183836 6180 183888 6186
rect 183836 6122 183888 6128
rect 185228 5982 185256 97922
rect 185320 16574 185348 99826
rect 185688 98122 185716 102037
rect 185676 98116 185728 98122
rect 185676 98058 185728 98064
rect 186148 97986 186176 102037
rect 186412 98048 186464 98054
rect 186412 97990 186464 97996
rect 186136 97980 186188 97986
rect 186136 97922 186188 97928
rect 186320 97980 186372 97986
rect 186320 97922 186372 97928
rect 185320 16546 186176 16574
rect 185216 5976 185268 5982
rect 185216 5918 185268 5924
rect 183652 4616 183704 4622
rect 183652 4558 183704 4564
rect 184940 3596 184992 3602
rect 184940 3538 184992 3544
rect 183572 3454 183784 3482
rect 183756 480 183784 3454
rect 184952 480 184980 3538
rect 186148 480 186176 16546
rect 186332 3806 186360 97922
rect 186424 6050 186452 97990
rect 186608 84194 186636 102037
rect 187068 97986 187096 102037
rect 187620 98054 187648 102037
rect 187608 98048 187660 98054
rect 187608 97990 187660 97996
rect 187056 97980 187108 97986
rect 188080 97968 188108 102037
rect 187056 97922 187108 97928
rect 187712 97940 188108 97968
rect 186516 84166 186636 84194
rect 186516 6730 186544 84166
rect 186504 6724 186556 6730
rect 186504 6666 186556 6672
rect 187712 6662 187740 97940
rect 188540 84194 188568 102037
rect 189092 100434 189120 102037
rect 188988 100428 189040 100434
rect 188988 100370 189040 100376
rect 189080 100428 189132 100434
rect 189080 100370 189132 100376
rect 189000 100314 189028 100370
rect 189000 100286 189120 100314
rect 187804 84166 188568 84194
rect 187804 7954 187832 84166
rect 187792 7948 187844 7954
rect 187792 7890 187844 7896
rect 187700 6656 187752 6662
rect 187700 6598 187752 6604
rect 186412 6044 186464 6050
rect 186412 5986 186464 5992
rect 187332 5432 187384 5438
rect 187332 5374 187384 5380
rect 186320 3800 186372 3806
rect 186320 3742 186372 3748
rect 187344 480 187372 5374
rect 188528 3528 188580 3534
rect 188528 3470 188580 3476
rect 188540 480 188568 3470
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189092 354 189120 100286
rect 189172 97980 189224 97986
rect 189172 97922 189224 97928
rect 189184 3738 189212 97922
rect 189552 84194 189580 102037
rect 190012 97986 190040 102037
rect 190000 97980 190052 97986
rect 190000 97922 190052 97928
rect 190460 97980 190512 97986
rect 190460 97922 190512 97928
rect 189276 84166 189580 84194
rect 189276 16574 189304 84166
rect 189276 16546 189396 16574
rect 189368 6594 189396 16546
rect 189356 6588 189408 6594
rect 189356 6530 189408 6536
rect 189172 3732 189224 3738
rect 189172 3674 189224 3680
rect 190472 3670 190500 97922
rect 190564 4486 190592 102037
rect 191024 84194 191052 102037
rect 191484 97986 191512 102037
rect 191472 97980 191524 97986
rect 191472 97922 191524 97928
rect 191840 97980 191892 97986
rect 191840 97922 191892 97928
rect 190656 84166 191052 84194
rect 190656 6526 190684 84166
rect 190644 6520 190696 6526
rect 190644 6462 190696 6468
rect 190828 5364 190880 5370
rect 190828 5306 190880 5312
rect 190552 4480 190604 4486
rect 190552 4422 190604 4428
rect 190460 3664 190512 3670
rect 190460 3606 190512 3612
rect 190840 480 190868 5306
rect 191852 3602 191880 97922
rect 191944 4690 191972 102037
rect 192496 84194 192524 102037
rect 192956 97986 192984 102037
rect 193220 100700 193272 100706
rect 193220 100642 193272 100648
rect 192944 97980 192996 97986
rect 192944 97922 192996 97928
rect 192036 84166 192524 84194
rect 192036 6254 192064 84166
rect 192024 6248 192076 6254
rect 192024 6190 192076 6196
rect 191932 4684 191984 4690
rect 191932 4626 191984 4632
rect 191840 3596 191892 3602
rect 191840 3538 191892 3544
rect 192024 3460 192076 3466
rect 192024 3402 192076 3408
rect 192036 480 192064 3402
rect 193232 480 193260 100642
rect 193416 98002 193444 102037
rect 193324 97974 193444 98002
rect 193324 4758 193352 97974
rect 193968 97866 193996 102037
rect 193416 97838 193996 97866
rect 193416 6458 193444 97838
rect 194428 84194 194456 102037
rect 194888 100706 194916 102037
rect 194876 100700 194928 100706
rect 194876 100642 194928 100648
rect 194600 97980 194652 97986
rect 194600 97922 194652 97928
rect 193508 84166 194456 84194
rect 193508 7886 193536 84166
rect 193496 7880 193548 7886
rect 193496 7822 193548 7828
rect 193404 6452 193456 6458
rect 193404 6394 193456 6400
rect 194416 5296 194468 5302
rect 194416 5238 194468 5244
rect 193312 4752 193364 4758
rect 193312 4694 193364 4700
rect 194428 480 194456 5238
rect 194612 3534 194640 97922
rect 195348 84194 195376 102037
rect 195900 97986 195928 102037
rect 196360 100570 196388 102037
rect 195980 100564 196032 100570
rect 195980 100506 196032 100512
rect 196348 100564 196400 100570
rect 196348 100506 196400 100512
rect 195888 97980 195940 97986
rect 195888 97922 195940 97928
rect 194704 84166 195376 84194
rect 194704 7818 194732 84166
rect 194692 7812 194744 7818
rect 194692 7754 194744 7760
rect 195612 4140 195664 4146
rect 195612 4082 195664 4088
rect 194600 3528 194652 3534
rect 194600 3470 194652 3476
rect 195624 480 195652 4082
rect 195992 3482 196020 100506
rect 196820 84194 196848 102037
rect 197372 98002 197400 102037
rect 197372 97974 197584 98002
rect 197452 97912 197504 97918
rect 197452 97854 197504 97860
rect 197360 97844 197412 97850
rect 197360 97786 197412 97792
rect 196084 84166 196848 84194
rect 196084 6390 196112 84166
rect 196072 6384 196124 6390
rect 196072 6326 196124 6332
rect 197372 5506 197400 97786
rect 197464 6322 197492 97854
rect 197556 7682 197584 97974
rect 197832 97850 197860 102037
rect 198292 97918 198320 102037
rect 198280 97912 198332 97918
rect 198280 97854 198332 97860
rect 197820 97844 197872 97850
rect 197820 97786 197872 97792
rect 197544 7676 197596 7682
rect 197544 7618 197596 7624
rect 197452 6316 197504 6322
rect 197452 6258 197504 6264
rect 197360 5500 197412 5506
rect 197360 5442 197412 5448
rect 197912 5228 197964 5234
rect 197912 5170 197964 5176
rect 195992 3454 196848 3482
rect 196820 480 196848 3454
rect 197924 480 197952 5170
rect 198752 3466 198780 102037
rect 199304 98002 199332 102037
rect 199384 99952 199436 99958
rect 199384 99894 199436 99900
rect 198844 97974 199332 98002
rect 198844 5438 198872 97974
rect 198924 97912 198976 97918
rect 198924 97854 198976 97860
rect 198936 7614 198964 97854
rect 198924 7608 198976 7614
rect 198924 7550 198976 7556
rect 198832 5432 198884 5438
rect 198832 5374 198884 5380
rect 199396 4146 199424 99894
rect 199764 97918 199792 102037
rect 200120 100496 200172 100502
rect 200120 100438 200172 100444
rect 199752 97912 199804 97918
rect 199752 97854 199804 97860
rect 200132 6914 200160 100438
rect 200224 97968 200252 102037
rect 200776 99754 200804 102037
rect 200764 99748 200816 99754
rect 200764 99690 200816 99696
rect 200224 97940 200344 97968
rect 200212 97844 200264 97850
rect 200212 97786 200264 97792
rect 200224 7342 200252 97786
rect 200212 7336 200264 7342
rect 200212 7278 200264 7284
rect 200316 7274 200344 97940
rect 201236 97850 201264 102037
rect 201696 97968 201724 102037
rect 202248 99890 202276 102037
rect 202236 99884 202288 99890
rect 202236 99826 202288 99832
rect 201512 97940 201724 97968
rect 201224 97844 201276 97850
rect 201224 97786 201276 97792
rect 201512 7750 201540 97940
rect 202708 84194 202736 102037
rect 202880 100156 202932 100162
rect 202880 100098 202932 100104
rect 201604 84166 202736 84194
rect 201604 8158 201632 84166
rect 201592 8152 201644 8158
rect 201592 8094 201644 8100
rect 201500 7744 201552 7750
rect 201500 7686 201552 7692
rect 200304 7268 200356 7274
rect 200304 7210 200356 7216
rect 200132 6886 200344 6914
rect 199384 4140 199436 4146
rect 199384 4082 199436 4088
rect 199108 4072 199160 4078
rect 199108 4014 199160 4020
rect 198740 3460 198792 3466
rect 198740 3402 198792 3408
rect 199120 480 199148 4014
rect 200316 480 200344 6886
rect 201500 5160 201552 5166
rect 201500 5102 201552 5108
rect 201512 480 201540 5102
rect 202696 4140 202748 4146
rect 202696 4082 202748 4088
rect 202708 480 202736 4082
rect 202892 490 202920 100098
rect 203064 98048 203116 98054
rect 203064 97990 203116 97996
rect 202972 97980 203024 97986
rect 202972 97922 203024 97928
rect 202984 5370 203012 97922
rect 203076 8090 203104 97990
rect 203168 9382 203196 102037
rect 203628 97986 203656 102037
rect 204180 98054 204208 102037
rect 204168 98048 204220 98054
rect 204168 97990 204220 97996
rect 203616 97980 203668 97986
rect 203616 97922 203668 97928
rect 204640 84194 204668 102037
rect 205100 99958 205128 102037
rect 205652 100162 205680 102037
rect 205640 100156 205692 100162
rect 205640 100098 205692 100104
rect 205088 99952 205140 99958
rect 205088 99894 205140 99900
rect 206112 84194 206140 102037
rect 206284 100632 206336 100638
rect 206284 100574 206336 100580
rect 204272 84166 204668 84194
rect 205652 84166 206140 84194
rect 203156 9376 203208 9382
rect 203156 9318 203208 9324
rect 204272 9314 204300 84166
rect 204260 9308 204312 9314
rect 204260 9250 204312 9256
rect 205652 9246 205680 84166
rect 205640 9240 205692 9246
rect 205640 9182 205692 9188
rect 203064 8084 203116 8090
rect 203064 8026 203116 8032
rect 202972 5364 203024 5370
rect 202972 5306 203024 5312
rect 205088 5092 205140 5098
rect 205088 5034 205140 5040
rect 189694 354 189806 480
rect 189092 326 189806 354
rect 189694 -960 189806 326
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 202892 462 203472 490
rect 205100 480 205128 5034
rect 206192 4004 206244 4010
rect 206192 3946 206244 3952
rect 206204 480 206232 3946
rect 206296 3398 206324 100574
rect 206572 100502 206600 102037
rect 206560 100496 206612 100502
rect 206560 100438 206612 100444
rect 207032 8022 207060 102037
rect 207584 84194 207612 102037
rect 208044 99822 208072 102037
rect 208504 101946 208532 102037
rect 208412 101918 208532 101946
rect 208412 100638 208440 101918
rect 208400 100632 208452 100638
rect 208400 100574 208452 100580
rect 209056 100178 209084 102037
rect 208964 100150 209084 100178
rect 208032 99816 208084 99822
rect 208032 99758 208084 99764
rect 208400 97980 208452 97986
rect 208400 97922 208452 97928
rect 207124 84166 207612 84194
rect 207124 9178 207152 84166
rect 207112 9172 207164 9178
rect 207112 9114 207164 9120
rect 207020 8016 207072 8022
rect 207020 7958 207072 7964
rect 208412 5302 208440 97922
rect 208964 84194 208992 100150
rect 209044 100020 209096 100026
rect 209044 99962 209096 99968
rect 208504 84166 208992 84194
rect 208504 9110 208532 84166
rect 208492 9104 208544 9110
rect 208492 9046 208544 9052
rect 208400 5296 208452 5302
rect 208400 5238 208452 5244
rect 208584 5024 208636 5030
rect 208584 4966 208636 4972
rect 206284 3392 206336 3398
rect 206284 3334 206336 3340
rect 207388 3392 207440 3398
rect 207388 3334 207440 3340
rect 207400 480 207428 3334
rect 208596 480 208624 4966
rect 209056 3194 209084 99962
rect 209516 97986 209544 102037
rect 209976 100026 210004 102037
rect 210436 100178 210464 102037
rect 210344 100150 210464 100178
rect 209964 100020 210016 100026
rect 209964 99962 210016 99968
rect 209504 97980 209556 97986
rect 209504 97922 209556 97928
rect 209780 97980 209832 97986
rect 209780 97922 209832 97928
rect 209792 5234 209820 97922
rect 210344 84194 210372 100150
rect 210424 100088 210476 100094
rect 210424 100030 210476 100036
rect 209884 84166 210372 84194
rect 209884 9042 209912 84166
rect 209872 9036 209924 9042
rect 209872 8978 209924 8984
rect 209780 5228 209832 5234
rect 209780 5170 209832 5176
rect 209780 4956 209832 4962
rect 209780 4898 209832 4904
rect 209044 3188 209096 3194
rect 209044 3130 209096 3136
rect 209792 480 209820 4898
rect 210436 3398 210464 100030
rect 210988 97986 211016 102037
rect 211448 100094 211476 102037
rect 211908 100450 211936 102037
rect 211724 100422 211936 100450
rect 211436 100088 211488 100094
rect 211436 100030 211488 100036
rect 210976 97980 211028 97986
rect 210976 97922 211028 97928
rect 211160 97980 211212 97986
rect 211160 97922 211212 97928
rect 211172 5098 211200 97922
rect 211724 84194 211752 100422
rect 211804 100292 211856 100298
rect 211804 100234 211856 100240
rect 211264 84166 211752 84194
rect 211264 8974 211292 84166
rect 211252 8968 211304 8974
rect 211252 8910 211304 8916
rect 211160 5092 211212 5098
rect 211160 5034 211212 5040
rect 210424 3392 210476 3398
rect 210424 3334 210476 3340
rect 211816 3194 211844 100234
rect 212460 97986 212488 102037
rect 212920 100298 212948 102037
rect 213380 100450 213408 102037
rect 213104 100422 213408 100450
rect 212908 100292 212960 100298
rect 212908 100234 212960 100240
rect 212448 97980 212500 97986
rect 212448 97922 212500 97928
rect 213104 84194 213132 100422
rect 213184 100360 213236 100366
rect 213184 100302 213236 100308
rect 212552 84166 213132 84194
rect 212552 8634 212580 84166
rect 212540 8628 212592 8634
rect 212540 8570 212592 8576
rect 212172 4888 212224 4894
rect 212172 4830 212224 4836
rect 210976 3188 211028 3194
rect 210976 3130 211028 3136
rect 211804 3188 211856 3194
rect 211804 3130 211856 3136
rect 210988 480 211016 3130
rect 212184 480 212212 4830
rect 213196 3058 213224 100302
rect 213932 5166 213960 102037
rect 214392 98002 214420 102037
rect 214024 97974 214420 98002
rect 214024 8702 214052 97974
rect 214852 84194 214880 102037
rect 214116 84166 214880 84194
rect 214116 10946 214144 84166
rect 214104 10940 214156 10946
rect 214104 10882 214156 10888
rect 214012 8696 214064 8702
rect 214012 8638 214064 8644
rect 213920 5160 213972 5166
rect 213920 5102 213972 5108
rect 215312 5030 215340 102037
rect 215864 98002 215892 102037
rect 215944 100224 215996 100230
rect 215944 100166 215996 100172
rect 215404 97974 215892 98002
rect 215404 8770 215432 97974
rect 215484 97912 215536 97918
rect 215484 97854 215536 97860
rect 215496 10878 215524 97854
rect 215484 10872 215536 10878
rect 215484 10814 215536 10820
rect 215392 8764 215444 8770
rect 215392 8706 215444 8712
rect 215668 6112 215720 6118
rect 215668 6054 215720 6060
rect 215300 5024 215352 5030
rect 215300 4966 215352 4972
rect 213368 3936 213420 3942
rect 213368 3878 213420 3884
rect 213184 3052 213236 3058
rect 213184 2994 213236 3000
rect 213380 480 213408 3878
rect 214472 3392 214524 3398
rect 214472 3334 214524 3340
rect 214484 480 214512 3334
rect 215680 480 215708 6054
rect 215956 4078 215984 100166
rect 216324 97918 216352 102037
rect 216784 98002 216812 102037
rect 216692 97974 216812 98002
rect 216312 97912 216364 97918
rect 216312 97854 216364 97860
rect 216692 4962 216720 97974
rect 216772 97912 216824 97918
rect 216772 97854 216824 97860
rect 216784 10810 216812 97854
rect 217336 84194 217364 102037
rect 217796 97918 217824 102037
rect 218256 98002 218284 102037
rect 218072 97974 218284 98002
rect 217784 97912 217836 97918
rect 217784 97854 217836 97860
rect 216876 84166 217364 84194
rect 216876 15910 216904 84166
rect 216864 15904 216916 15910
rect 216864 15846 216916 15852
rect 216772 10804 216824 10810
rect 216772 10746 216824 10752
rect 218072 6914 218100 97974
rect 218152 97912 218204 97918
rect 218152 97854 218204 97860
rect 218164 10674 218192 97854
rect 218716 84194 218744 102037
rect 219268 97918 219296 102037
rect 219728 98002 219756 102037
rect 220188 100586 220216 102037
rect 219452 97974 219756 98002
rect 220004 100558 220216 100586
rect 219256 97912 219308 97918
rect 219256 97854 219308 97860
rect 218256 84166 218744 84194
rect 218256 10742 218284 84166
rect 218244 10736 218296 10742
rect 218244 10678 218296 10684
rect 218152 10668 218204 10674
rect 218152 10610 218204 10616
rect 218072 6886 218192 6914
rect 218060 6044 218112 6050
rect 218060 5986 218112 5992
rect 216772 5976 216824 5982
rect 216772 5918 216824 5924
rect 216680 4956 216732 4962
rect 216680 4898 216732 4904
rect 215944 4072 215996 4078
rect 215944 4014 215996 4020
rect 216784 4010 216812 5918
rect 216864 4820 216916 4826
rect 216864 4762 216916 4768
rect 216772 4004 216824 4010
rect 216772 3946 216824 3952
rect 216876 480 216904 4762
rect 218072 3942 218100 5986
rect 218164 4894 218192 6886
rect 218152 4888 218204 4894
rect 219452 4865 219480 97974
rect 220004 97900 220032 100558
rect 220084 100428 220136 100434
rect 220084 100370 220136 100376
rect 219544 97872 220032 97900
rect 219544 10606 219572 97872
rect 219624 97776 219676 97782
rect 219624 97718 219676 97724
rect 219532 10600 219584 10606
rect 219532 10542 219584 10548
rect 219636 10538 219664 97718
rect 219624 10532 219676 10538
rect 219624 10474 219676 10480
rect 218152 4830 218204 4836
rect 219438 4856 219494 4865
rect 219438 4791 219494 4800
rect 219256 4548 219308 4554
rect 219256 4490 219308 4496
rect 218060 3936 218112 3942
rect 218060 3878 218112 3884
rect 218060 3188 218112 3194
rect 218060 3130 218112 3136
rect 218072 480 218100 3130
rect 219268 480 219296 4490
rect 220096 4146 220124 100370
rect 220740 97782 220768 102037
rect 221200 98002 221228 102037
rect 220832 97974 221228 98002
rect 220728 97776 220780 97782
rect 220728 97718 220780 97724
rect 220832 4826 220860 97974
rect 220912 97912 220964 97918
rect 220912 97854 220964 97860
rect 220924 10334 220952 97854
rect 221660 84194 221688 102037
rect 222120 97918 222148 102037
rect 222672 100366 222700 102037
rect 222660 100360 222712 100366
rect 222660 100302 222712 100308
rect 222108 97912 222160 97918
rect 222108 97854 222160 97860
rect 223132 84194 223160 102037
rect 221016 84166 221688 84194
rect 222212 84166 223160 84194
rect 221016 10470 221044 84166
rect 221004 10464 221056 10470
rect 221004 10406 221056 10412
rect 222212 10402 222240 84166
rect 222200 10396 222252 10402
rect 222200 10338 222252 10344
rect 220912 10328 220964 10334
rect 220912 10270 220964 10276
rect 223592 9926 223620 102037
rect 224144 100434 224172 102037
rect 224224 100700 224276 100706
rect 224224 100642 224276 100648
rect 224132 100428 224184 100434
rect 224132 100370 224184 100376
rect 223580 9920 223632 9926
rect 223580 9862 223632 9868
rect 222752 6180 222804 6186
rect 222752 6122 222804 6128
rect 220820 4820 220872 4826
rect 220820 4762 220872 4768
rect 221740 4616 221792 4622
rect 221740 4558 221792 4564
rect 220084 4140 220136 4146
rect 220084 4082 220136 4088
rect 220544 4140 220596 4146
rect 220544 4082 220596 4088
rect 220556 3874 220584 4082
rect 220452 3868 220504 3874
rect 220452 3810 220504 3816
rect 220544 3868 220596 3874
rect 220544 3810 220596 3816
rect 220464 480 220492 3810
rect 221556 3052 221608 3058
rect 221556 2994 221608 3000
rect 221568 480 221596 2994
rect 221752 2854 221780 4558
rect 222476 4480 222528 4486
rect 222476 4422 222528 4428
rect 222488 3262 222516 4422
rect 222476 3256 222528 3262
rect 222476 3198 222528 3204
rect 221740 2848 221792 2854
rect 221740 2790 221792 2796
rect 222764 480 222792 6122
rect 224236 3330 224264 100642
rect 224604 100230 224632 102037
rect 224592 100224 224644 100230
rect 224592 100166 224644 100172
rect 224960 97980 225012 97986
rect 224960 97922 225012 97928
rect 224972 6186 225000 97922
rect 225064 9994 225092 102037
rect 225512 100564 225564 100570
rect 225512 100506 225564 100512
rect 225144 98048 225196 98054
rect 225144 97990 225196 97996
rect 225156 10062 225184 97990
rect 225524 93854 225552 100506
rect 225616 97986 225644 102037
rect 226076 98054 226104 102037
rect 226064 98048 226116 98054
rect 226064 97990 226116 97996
rect 226432 98048 226484 98054
rect 226432 97990 226484 97996
rect 225604 97980 225656 97986
rect 225604 97922 225656 97928
rect 226340 97980 226392 97986
rect 226340 97922 226392 97928
rect 225524 93826 225644 93854
rect 225144 10056 225196 10062
rect 225144 9998 225196 10004
rect 225052 9988 225104 9994
rect 225052 9930 225104 9936
rect 224960 6180 225012 6186
rect 224960 6122 225012 6128
rect 225144 4072 225196 4078
rect 225144 4014 225196 4020
rect 224224 3324 224276 3330
rect 224224 3266 224276 3272
rect 223948 2848 224000 2854
rect 223948 2790 224000 2796
rect 223960 480 223988 2790
rect 225156 480 225184 4014
rect 225616 3398 225644 93826
rect 226352 5914 226380 97922
rect 226444 10130 226472 97990
rect 226536 11558 226564 102037
rect 226892 99748 226944 99754
rect 226892 99690 226944 99696
rect 226904 93854 226932 99690
rect 226996 97986 227024 102037
rect 227548 98054 227576 102037
rect 227536 98048 227588 98054
rect 228008 98002 228036 102037
rect 227536 97990 227588 97996
rect 226984 97980 227036 97986
rect 226984 97922 227036 97928
rect 227720 97980 227772 97986
rect 227720 97922 227772 97928
rect 227824 97974 228036 98002
rect 228468 97986 228496 102037
rect 228456 97980 228508 97986
rect 226904 93826 227024 93854
rect 226524 11552 226576 11558
rect 226524 11494 226576 11500
rect 226432 10124 226484 10130
rect 226432 10066 226484 10072
rect 226432 6792 226484 6798
rect 226432 6734 226484 6740
rect 226340 5908 226392 5914
rect 226340 5850 226392 5856
rect 226444 3482 226472 6734
rect 226996 4078 227024 93826
rect 227536 6860 227588 6866
rect 227536 6802 227588 6808
rect 226984 4072 227036 4078
rect 226984 4014 227036 4020
rect 226352 3454 226472 3482
rect 225604 3392 225656 3398
rect 225604 3334 225656 3340
rect 226352 480 226380 3454
rect 227548 480 227576 6802
rect 227732 5982 227760 97922
rect 227824 14278 227852 97974
rect 228456 97922 228508 97928
rect 229020 84194 229048 102037
rect 229100 98116 229152 98122
rect 229100 98058 229152 98064
rect 227916 84166 229048 84194
rect 227916 18426 227944 84166
rect 227904 18420 227956 18426
rect 227904 18362 227956 18368
rect 227812 14272 227864 14278
rect 227812 14214 227864 14220
rect 229112 6050 229140 98058
rect 229480 98002 229508 102037
rect 229744 99884 229796 99890
rect 229744 99826 229796 99832
rect 229204 97974 229508 98002
rect 229204 15706 229232 97974
rect 229284 97912 229336 97918
rect 229284 97854 229336 97860
rect 229296 18494 229324 97854
rect 229284 18488 229336 18494
rect 229284 18430 229336 18436
rect 229192 15700 229244 15706
rect 229192 15642 229244 15648
rect 229100 6044 229152 6050
rect 229100 5986 229152 5992
rect 227720 5976 227772 5982
rect 227720 5918 227772 5924
rect 229756 4010 229784 99826
rect 229940 98122 229968 102037
rect 229928 98116 229980 98122
rect 229928 98058 229980 98064
rect 230400 97918 230428 102037
rect 230480 97980 230532 97986
rect 230480 97922 230532 97928
rect 230388 97912 230440 97918
rect 230388 97854 230440 97860
rect 229836 6724 229888 6730
rect 229836 6666 229888 6672
rect 228732 4004 228784 4010
rect 228732 3946 228784 3952
rect 229744 4004 229796 4010
rect 229744 3946 229796 3952
rect 228744 480 228772 3946
rect 229848 480 229876 6666
rect 230492 6118 230520 97922
rect 230952 84194 230980 102037
rect 231412 97986 231440 102037
rect 231400 97980 231452 97986
rect 231400 97922 231452 97928
rect 231872 97918 231900 102037
rect 232424 98002 232452 102037
rect 232504 99952 232556 99958
rect 232504 99894 232556 99900
rect 231964 97974 232452 98002
rect 231860 97912 231912 97918
rect 231860 97854 231912 97860
rect 231860 97776 231912 97782
rect 231860 97718 231912 97724
rect 230584 84166 230980 84194
rect 230584 15774 230612 84166
rect 230572 15768 230624 15774
rect 230572 15710 230624 15716
rect 231872 6866 231900 97718
rect 231964 15842 231992 97974
rect 232044 97912 232096 97918
rect 232044 97854 232096 97860
rect 232056 19786 232084 97854
rect 232044 19780 232096 19786
rect 232044 19722 232096 19728
rect 231952 15836 232004 15842
rect 231952 15778 232004 15784
rect 231860 6860 231912 6866
rect 231860 6802 231912 6808
rect 230480 6112 230532 6118
rect 230480 6054 230532 6060
rect 232516 4146 232544 99894
rect 232884 97782 232912 102037
rect 233240 97980 233292 97986
rect 233240 97922 233292 97928
rect 232872 97776 232924 97782
rect 232872 97718 232924 97724
rect 233252 6798 233280 97922
rect 233344 11626 233372 102037
rect 233804 84194 233832 102037
rect 233884 99816 233936 99822
rect 233884 99758 233936 99764
rect 233436 84166 233832 84194
rect 233436 16590 233464 84166
rect 233424 16584 233476 16590
rect 233424 16526 233476 16532
rect 233332 11620 233384 11626
rect 233332 11562 233384 11568
rect 233240 6792 233292 6798
rect 233240 6734 233292 6740
rect 233424 6656 233476 6662
rect 233424 6598 233476 6604
rect 232504 4140 232556 4146
rect 232504 4082 232556 4088
rect 232228 3936 232280 3942
rect 232228 3878 232280 3884
rect 231032 3800 231084 3806
rect 231032 3742 231084 3748
rect 231044 480 231072 3742
rect 232240 480 232268 3878
rect 233436 480 233464 6598
rect 233896 3806 233924 99758
rect 234356 97986 234384 102037
rect 234816 98002 234844 102037
rect 235276 98002 235304 102037
rect 235356 100496 235408 100502
rect 235356 100438 235408 100444
rect 234344 97980 234396 97986
rect 234344 97922 234396 97928
rect 234620 97980 234672 97986
rect 234620 97922 234672 97928
rect 234724 97974 234844 98002
rect 235184 97974 235304 98002
rect 234632 6730 234660 97922
rect 234724 11694 234752 97974
rect 235184 84194 235212 97974
rect 235368 84194 235396 100438
rect 235828 97986 235856 102037
rect 236288 99634 236316 102037
rect 236104 99606 236316 99634
rect 235816 97980 235868 97986
rect 235816 97922 235868 97928
rect 234816 84166 235212 84194
rect 235276 84166 235396 84194
rect 234816 19854 234844 84166
rect 234804 19848 234856 19854
rect 234804 19790 234856 19796
rect 234712 11688 234764 11694
rect 234712 11630 234764 11636
rect 234712 7948 234764 7954
rect 234712 7890 234764 7896
rect 234620 6724 234672 6730
rect 234620 6666 234672 6672
rect 233884 3800 233936 3806
rect 233884 3742 233936 3748
rect 234724 3482 234752 7890
rect 235276 3942 235304 84166
rect 236104 12442 236132 99606
rect 236748 98002 236776 102037
rect 236196 97974 236776 98002
rect 236196 21214 236224 97974
rect 237300 84194 237328 102037
rect 237760 98002 237788 102037
rect 238220 100722 238248 102037
rect 236288 84166 237328 84194
rect 237392 97974 237788 98002
rect 237944 100694 238248 100722
rect 236184 21208 236236 21214
rect 236184 21150 236236 21156
rect 236092 12436 236144 12442
rect 236092 12378 236144 12384
rect 236288 6225 236316 84166
rect 237392 12374 237420 97974
rect 237472 97912 237524 97918
rect 237472 97854 237524 97860
rect 237484 17066 237512 97854
rect 237944 84194 237972 100694
rect 238024 100632 238076 100638
rect 238024 100574 238076 100580
rect 237576 84166 237972 84194
rect 237576 21282 237604 84166
rect 237564 21276 237616 21282
rect 237564 21218 237616 21224
rect 237472 17060 237524 17066
rect 237472 17002 237524 17008
rect 237380 12368 237432 12374
rect 237380 12310 237432 12316
rect 237380 8152 237432 8158
rect 237380 8094 237432 8100
rect 237012 6588 237064 6594
rect 237012 6530 237064 6536
rect 236274 6216 236330 6225
rect 236274 6151 236330 6160
rect 235264 3936 235316 3942
rect 235264 3878 235316 3884
rect 235816 3868 235868 3874
rect 235816 3810 235868 3816
rect 234632 3454 234752 3482
rect 234632 480 234660 3454
rect 235828 480 235856 3810
rect 237024 480 237052 6530
rect 237392 3874 237420 8094
rect 238036 5778 238064 100574
rect 238680 97918 238708 102037
rect 239232 97968 239260 102037
rect 238772 97940 239260 97968
rect 238668 97912 238720 97918
rect 238668 97854 238720 97860
rect 238772 12306 238800 97940
rect 239692 84194 239720 102037
rect 240152 97968 240180 102037
rect 240152 97940 240272 97968
rect 240140 97844 240192 97850
rect 240140 97786 240192 97792
rect 238864 84166 239720 84194
rect 238864 21350 238892 84166
rect 238852 21344 238904 21350
rect 238852 21286 238904 21292
rect 238760 12300 238812 12306
rect 238760 12242 238812 12248
rect 240152 12238 240180 97786
rect 240244 17134 240272 97940
rect 240704 97850 240732 102037
rect 240692 97844 240744 97850
rect 240692 97786 240744 97792
rect 241164 84194 241192 102037
rect 241520 97980 241572 97986
rect 241520 97922 241572 97928
rect 240336 84166 241192 84194
rect 240336 22098 240364 84166
rect 240324 22092 240376 22098
rect 240324 22034 240376 22040
rect 240232 17128 240284 17134
rect 240232 17070 240284 17076
rect 240140 12232 240192 12238
rect 240140 12174 240192 12180
rect 241532 12170 241560 97922
rect 241624 17202 241652 102037
rect 241704 101788 241756 101794
rect 241704 101730 241756 101736
rect 241716 22030 241744 101730
rect 242084 97986 242112 102037
rect 242636 101794 242664 102037
rect 242624 101788 242676 101794
rect 242624 101730 242676 101736
rect 242164 100360 242216 100366
rect 242164 100302 242216 100308
rect 242072 97980 242124 97986
rect 242072 97922 242124 97928
rect 241704 22024 241756 22030
rect 241704 21966 241756 21972
rect 241612 17196 241664 17202
rect 241612 17138 241664 17144
rect 241520 12164 241572 12170
rect 241520 12106 241572 12112
rect 240140 8084 240192 8090
rect 240140 8026 240192 8032
rect 238024 5772 238076 5778
rect 238024 5714 238076 5720
rect 237380 3868 237432 3874
rect 237380 3810 237432 3816
rect 240152 3738 240180 8026
rect 240508 6520 240560 6526
rect 240508 6462 240560 6468
rect 238116 3732 238168 3738
rect 238116 3674 238168 3680
rect 240140 3732 240192 3738
rect 240140 3674 240192 3680
rect 238128 480 238156 3674
rect 239312 3256 239364 3262
rect 239312 3198 239364 3204
rect 239324 480 239352 3198
rect 240520 480 240548 6462
rect 242176 4554 242204 100302
rect 242900 97980 242952 97986
rect 243096 97968 243124 102037
rect 243360 100428 243412 100434
rect 243360 100370 243412 100376
rect 242900 97922 242952 97928
rect 243004 97940 243124 97968
rect 242912 12102 242940 97922
rect 243004 17950 243032 97940
rect 243084 97844 243136 97850
rect 243084 97786 243136 97792
rect 243096 21962 243124 97786
rect 243372 97730 243400 100370
rect 243556 97986 243584 102037
rect 243636 100292 243688 100298
rect 243636 100234 243688 100240
rect 243544 97980 243596 97986
rect 243544 97922 243596 97928
rect 243372 97702 243584 97730
rect 243084 21956 243136 21962
rect 243084 21898 243136 21904
rect 242992 17944 243044 17950
rect 242992 17886 243044 17892
rect 242900 12096 242952 12102
rect 242900 12038 242952 12044
rect 242900 4684 242952 4690
rect 242900 4626 242952 4632
rect 242164 4548 242216 4554
rect 242164 4490 242216 4496
rect 241704 3664 241756 3670
rect 241704 3606 241756 3612
rect 241716 480 241744 3606
rect 242912 480 242940 4626
rect 243556 4622 243584 97702
rect 243648 5846 243676 100234
rect 244108 97850 244136 102037
rect 244280 97980 244332 97986
rect 244568 97968 244596 102037
rect 245028 97986 245056 102037
rect 244280 97922 244332 97928
rect 244384 97940 244596 97968
rect 245016 97980 245068 97986
rect 244096 97844 244148 97850
rect 244096 97786 244148 97792
rect 244292 12034 244320 97922
rect 244384 17882 244412 97940
rect 245016 97922 245068 97928
rect 245580 84194 245608 102037
rect 246040 97968 246068 102037
rect 246500 100314 246528 102037
rect 244476 84166 245608 84194
rect 245672 97940 246068 97968
rect 246224 100286 246528 100314
rect 244476 21894 244504 84166
rect 244464 21888 244516 21894
rect 244464 21830 244516 21836
rect 244372 17876 244424 17882
rect 244372 17818 244424 17824
rect 244280 12028 244332 12034
rect 244280 11970 244332 11976
rect 245672 7410 245700 97940
rect 246224 97900 246252 100286
rect 246304 100224 246356 100230
rect 246304 100166 246356 100172
rect 245764 97872 246252 97900
rect 245764 11966 245792 97872
rect 245844 97776 245896 97782
rect 245844 97718 245896 97724
rect 245856 21826 245884 97718
rect 245844 21820 245896 21826
rect 245844 21762 245896 21768
rect 245752 11960 245804 11966
rect 245752 11902 245804 11908
rect 245660 7404 245712 7410
rect 245660 7346 245712 7352
rect 246316 6254 246344 100166
rect 246960 97782 246988 102037
rect 247512 97968 247540 102037
rect 247972 100314 248000 102037
rect 248432 100722 248460 102037
rect 248432 100694 248644 100722
rect 247052 97940 247540 97968
rect 247604 100286 248000 100314
rect 246948 97776 247000 97782
rect 246948 97718 247000 97724
rect 247052 7478 247080 97940
rect 247604 84194 247632 100286
rect 247684 100156 247736 100162
rect 247684 100098 247736 100104
rect 247144 84166 247632 84194
rect 247144 11898 247172 84166
rect 247132 11892 247184 11898
rect 247132 11834 247184 11840
rect 247040 7472 247092 7478
rect 247040 7414 247092 7420
rect 247592 6452 247644 6458
rect 247592 6394 247644 6400
rect 244096 6248 244148 6254
rect 244096 6190 244148 6196
rect 246304 6248 246356 6254
rect 246304 6190 246356 6196
rect 243636 5840 243688 5846
rect 243636 5782 243688 5788
rect 243544 4616 243596 4622
rect 243544 4558 243596 4564
rect 243452 4208 243504 4214
rect 243452 4150 243504 4156
rect 243464 3874 243492 4150
rect 243636 4140 243688 4146
rect 243636 4082 243688 4088
rect 243648 3942 243676 4082
rect 243636 3936 243688 3942
rect 243636 3878 243688 3884
rect 243452 3868 243504 3874
rect 243452 3810 243504 3816
rect 244108 480 244136 6190
rect 246396 4752 246448 4758
rect 246396 4694 246448 4700
rect 245200 3596 245252 3602
rect 245200 3538 245252 3544
rect 245212 480 245240 3538
rect 246408 480 246436 4694
rect 247604 480 247632 6394
rect 247696 3602 247724 100098
rect 248328 99476 248380 99482
rect 248328 99418 248380 99424
rect 248340 99090 248368 99418
rect 248340 99062 248460 99090
rect 248432 7546 248460 99062
rect 248512 97980 248564 97986
rect 248512 97922 248564 97928
rect 248524 11830 248552 97922
rect 248616 21758 248644 100694
rect 248984 99482 249012 102037
rect 248972 99476 249024 99482
rect 248972 99418 249024 99424
rect 249444 97986 249472 102037
rect 249800 98252 249852 98258
rect 249800 98194 249852 98200
rect 249432 97980 249484 97986
rect 249432 97922 249484 97928
rect 248604 21752 248656 21758
rect 248604 21694 248656 21700
rect 248512 11824 248564 11830
rect 248512 11766 248564 11772
rect 249812 8294 249840 98194
rect 249904 98002 249932 102037
rect 250364 98258 250392 102037
rect 250352 98252 250404 98258
rect 250352 98194 250404 98200
rect 249904 97974 250024 98002
rect 249892 97912 249944 97918
rect 249892 97854 249944 97860
rect 249904 11762 249932 97854
rect 249996 21690 250024 97974
rect 250916 97918 250944 102037
rect 251272 98048 251324 98054
rect 251272 97990 251324 97996
rect 251180 97980 251232 97986
rect 251180 97922 251232 97928
rect 250904 97912 250956 97918
rect 250904 97854 250956 97860
rect 249984 21684 250036 21690
rect 249984 21626 250036 21632
rect 249892 11756 249944 11762
rect 249892 11698 249944 11704
rect 249800 8288 249852 8294
rect 249800 8230 249852 8236
rect 251192 8226 251220 97922
rect 251284 19922 251312 97990
rect 251376 21622 251404 102037
rect 251836 97986 251864 102037
rect 252388 98054 252416 102037
rect 252848 100366 252876 102037
rect 252836 100360 252888 100366
rect 252836 100302 252888 100308
rect 252376 98048 252428 98054
rect 253308 98002 253336 102037
rect 252376 97990 252428 97996
rect 251824 97980 251876 97986
rect 251824 97922 251876 97928
rect 252572 97974 253336 98002
rect 251364 21616 251416 21622
rect 251364 21558 251416 21564
rect 251272 19916 251324 19922
rect 251272 19858 251324 19864
rect 251180 8220 251232 8226
rect 251180 8162 251232 8168
rect 252572 8158 252600 97974
rect 253768 84194 253796 102037
rect 254032 98048 254084 98054
rect 254032 97990 254084 97996
rect 253940 97980 253992 97986
rect 253940 97922 253992 97928
rect 252664 84166 253796 84194
rect 252664 20602 252692 84166
rect 252652 20596 252704 20602
rect 252652 20538 252704 20544
rect 252560 8152 252612 8158
rect 252560 8094 252612 8100
rect 253952 8090 253980 97922
rect 254044 20534 254072 97990
rect 254320 84194 254348 102037
rect 254780 97986 254808 102037
rect 255240 98054 255268 102037
rect 255792 100298 255820 102037
rect 255780 100292 255832 100298
rect 255780 100234 255832 100240
rect 255228 98048 255280 98054
rect 255228 97990 255280 97996
rect 254768 97980 254820 97986
rect 254768 97922 254820 97928
rect 256252 84194 256280 102037
rect 256712 98002 256740 102037
rect 256712 97974 256832 98002
rect 256700 97912 256752 97918
rect 256700 97854 256752 97860
rect 254136 84166 254348 84194
rect 255332 84166 256280 84194
rect 254136 23186 254164 84166
rect 254124 23180 254176 23186
rect 254124 23122 254176 23128
rect 254032 20528 254084 20534
rect 254032 20470 254084 20476
rect 253940 8084 253992 8090
rect 253940 8026 253992 8032
rect 255332 8022 255360 84166
rect 249800 8016 249852 8022
rect 249800 7958 249852 7964
rect 255320 8016 255372 8022
rect 255320 7958 255372 7964
rect 248788 7880 248840 7886
rect 248788 7822 248840 7828
rect 248420 7540 248472 7546
rect 248420 7482 248472 7488
rect 247684 3596 247736 3602
rect 247684 3538 247736 3544
rect 248800 480 248828 7822
rect 249812 3670 249840 7958
rect 256712 7954 256740 97854
rect 256804 20466 256832 97974
rect 257264 84194 257292 102037
rect 257344 100088 257396 100094
rect 257344 100030 257396 100036
rect 256896 84166 257292 84194
rect 256896 23118 256924 84166
rect 256884 23112 256936 23118
rect 256884 23054 256936 23060
rect 256792 20460 256844 20466
rect 256792 20402 256844 20408
rect 256700 7948 256752 7954
rect 256700 7890 256752 7896
rect 251180 7812 251232 7818
rect 251180 7754 251232 7760
rect 249800 3664 249852 3670
rect 249800 3606 249852 3612
rect 249984 3324 250036 3330
rect 249984 3266 250036 3272
rect 249996 480 250024 3266
rect 251192 480 251220 7754
rect 255872 7676 255924 7682
rect 255872 7618 255924 7624
rect 254676 6384 254728 6390
rect 254676 6326 254728 6332
rect 252376 3528 252428 3534
rect 252376 3470 252428 3476
rect 252388 480 252416 3470
rect 253480 3392 253532 3398
rect 253480 3334 253532 3340
rect 253492 480 253520 3334
rect 254688 480 254716 6326
rect 255884 480 255912 7618
rect 257356 5506 257384 100030
rect 257436 100020 257488 100026
rect 257436 99962 257488 99968
rect 257068 5500 257120 5506
rect 257068 5442 257120 5448
rect 257344 5500 257396 5506
rect 257344 5442 257396 5448
rect 257080 480 257108 5442
rect 257448 4758 257476 99962
rect 257724 97918 257752 102037
rect 258080 97980 258132 97986
rect 258080 97922 258132 97928
rect 257712 97912 257764 97918
rect 257712 97854 257764 97860
rect 258092 7886 258120 97922
rect 258184 20398 258212 102037
rect 258644 100230 258672 102037
rect 258632 100224 258684 100230
rect 258632 100166 258684 100172
rect 259196 97986 259224 102037
rect 259184 97980 259236 97986
rect 259184 97922 259236 97928
rect 259460 97980 259512 97986
rect 259656 97968 259684 102037
rect 259460 97922 259512 97928
rect 259564 97940 259684 97968
rect 258172 20392 258224 20398
rect 258172 20334 258224 20340
rect 258080 7880 258132 7886
rect 258080 7822 258132 7828
rect 259472 7818 259500 97922
rect 259564 12918 259592 97940
rect 260116 84194 260144 102037
rect 260668 97986 260696 102037
rect 260656 97980 260708 97986
rect 260656 97922 260708 97928
rect 260840 97980 260892 97986
rect 260840 97922 260892 97928
rect 259656 84166 260144 84194
rect 259656 23050 259684 84166
rect 259644 23044 259696 23050
rect 259644 22986 259696 22992
rect 259552 12912 259604 12918
rect 259552 12854 259604 12860
rect 259460 7812 259512 7818
rect 259460 7754 259512 7760
rect 260852 7750 260880 97922
rect 261128 84194 261156 102037
rect 261588 100162 261616 102037
rect 261576 100156 261628 100162
rect 261576 100098 261628 100104
rect 262048 97986 262076 102037
rect 262036 97980 262088 97986
rect 262036 97922 262088 97928
rect 262220 97980 262272 97986
rect 262600 97968 262628 102037
rect 262220 97922 262272 97928
rect 262324 97940 262628 97968
rect 260944 84166 261156 84194
rect 260944 12986 260972 84166
rect 260932 12980 260984 12986
rect 260932 12922 260984 12928
rect 258080 7744 258132 7750
rect 258080 7686 258132 7692
rect 260840 7744 260892 7750
rect 260840 7686 260892 7692
rect 257436 4752 257488 4758
rect 257436 4694 257488 4700
rect 258092 3534 258120 7686
rect 262232 7682 262260 97922
rect 262324 13054 262352 97940
rect 263060 84194 263088 102037
rect 263520 97986 263548 102037
rect 263508 97980 263560 97986
rect 263508 97922 263560 97928
rect 264072 84194 264100 102037
rect 264532 100502 264560 102037
rect 264520 100496 264572 100502
rect 264520 100438 264572 100444
rect 262416 84166 263088 84194
rect 263612 84166 264100 84194
rect 262416 22982 262444 84166
rect 262404 22976 262456 22982
rect 262404 22918 262456 22924
rect 263612 13802 263640 84166
rect 263600 13796 263652 13802
rect 263600 13738 263652 13744
rect 262312 13048 262364 13054
rect 262312 12990 262364 12996
rect 262220 7676 262272 7682
rect 262220 7618 262272 7624
rect 264992 7614 265020 102037
rect 265452 97968 265480 102037
rect 265084 97940 265480 97968
rect 265084 13734 265112 97940
rect 266004 84194 266032 102037
rect 266360 97980 266412 97986
rect 266360 97922 266412 97928
rect 265176 84166 266032 84194
rect 265176 22914 265204 84166
rect 265164 22908 265216 22914
rect 265164 22850 265216 22856
rect 265072 13728 265124 13734
rect 265072 13670 265124 13676
rect 266372 13666 266400 97922
rect 266464 18562 266492 102037
rect 266924 97986 266952 102037
rect 267476 100094 267504 102037
rect 267464 100088 267516 100094
rect 267464 100030 267516 100036
rect 267936 98002 267964 102037
rect 266912 97980 266964 97986
rect 266912 97922 266964 97928
rect 267740 97980 267792 97986
rect 267740 97922 267792 97928
rect 267844 97974 267964 98002
rect 268396 97986 268424 102037
rect 268384 97980 268436 97986
rect 266452 18556 266504 18562
rect 266452 18498 266504 18504
rect 266360 13660 266412 13666
rect 266360 13602 266412 13608
rect 267752 13598 267780 97922
rect 267844 19310 267872 97974
rect 268384 97922 268436 97928
rect 268948 84194 268976 102037
rect 269120 97980 269172 97986
rect 269120 97922 269172 97928
rect 267936 84166 268976 84194
rect 267936 22846 267964 84166
rect 267924 22840 267976 22846
rect 267924 22782 267976 22788
rect 267832 19304 267884 19310
rect 267832 19246 267884 19252
rect 267740 13592 267792 13598
rect 267740 13534 267792 13540
rect 269132 13530 269160 97922
rect 269408 84194 269436 102037
rect 269868 97986 269896 102037
rect 270328 100026 270356 102037
rect 270316 100020 270368 100026
rect 270316 99962 270368 99968
rect 270880 98002 270908 102037
rect 269856 97980 269908 97986
rect 269856 97922 269908 97928
rect 270500 97980 270552 97986
rect 270500 97922 270552 97928
rect 270604 97974 270908 98002
rect 271340 97986 271368 102037
rect 271328 97980 271380 97986
rect 269224 84166 269436 84194
rect 269224 19242 269252 84166
rect 269212 19236 269264 19242
rect 269212 19178 269264 19184
rect 269120 13524 269172 13530
rect 269120 13466 269172 13472
rect 270512 13462 270540 97922
rect 270604 19174 270632 97974
rect 271328 97922 271380 97928
rect 271800 84194 271828 102037
rect 271880 97980 271932 97986
rect 271880 97922 271932 97928
rect 270696 84166 271828 84194
rect 270696 22778 270724 84166
rect 270684 22772 270736 22778
rect 270684 22714 270736 22720
rect 270592 19168 270644 19174
rect 270592 19110 270644 19116
rect 270500 13456 270552 13462
rect 270500 13398 270552 13404
rect 271892 13394 271920 97922
rect 272352 84194 272380 102037
rect 272812 97986 272840 102037
rect 272800 97980 272852 97986
rect 272800 97922 272852 97928
rect 271984 84166 272380 84194
rect 271984 19106 272012 84166
rect 271972 19100 272024 19106
rect 271972 19042 272024 19048
rect 271880 13388 271932 13394
rect 271880 13330 271932 13336
rect 270040 9376 270092 9382
rect 270040 9318 270092 9324
rect 261760 7608 261812 7614
rect 261760 7550 261812 7556
rect 264980 7608 265032 7614
rect 264980 7550 265032 7556
rect 258264 6316 258316 6322
rect 258264 6258 258316 6264
rect 258080 3528 258132 3534
rect 258080 3470 258132 3476
rect 258276 480 258304 6258
rect 260656 5432 260708 5438
rect 260656 5374 260708 5380
rect 259460 3460 259512 3466
rect 259460 3402 259512 3408
rect 259472 480 259500 3402
rect 260668 480 260696 5374
rect 261772 480 261800 7550
rect 265348 7336 265400 7342
rect 265348 7278 265400 7284
rect 262956 7268 263008 7274
rect 262956 7210 263008 7216
rect 262968 480 262996 7210
rect 264152 4072 264204 4078
rect 264152 4014 264204 4020
rect 264164 480 264192 4014
rect 265360 480 265388 7278
rect 268844 4140 268896 4146
rect 268844 4082 268896 4088
rect 267740 4004 267792 4010
rect 267740 3946 267792 3952
rect 266544 3528 266596 3534
rect 266544 3470 266596 3476
rect 266556 480 266584 3470
rect 267752 480 267780 3946
rect 268856 480 268884 4082
rect 270052 480 270080 9318
rect 271236 5364 271288 5370
rect 271236 5306 271288 5312
rect 271248 480 271276 5306
rect 272432 3732 272484 3738
rect 272432 3674 272484 3680
rect 272444 480 272472 3674
rect 273272 3262 273300 102037
rect 273732 98002 273760 102037
rect 273364 97974 273760 98002
rect 273364 8838 273392 97974
rect 274284 84194 274312 102037
rect 274744 98002 274772 102037
rect 273456 84166 274312 84194
rect 274652 97974 274772 98002
rect 273456 13326 273484 84166
rect 273444 13320 273496 13326
rect 273444 13262 273496 13268
rect 273628 9308 273680 9314
rect 273628 9250 273680 9256
rect 273352 8832 273404 8838
rect 273352 8774 273404 8780
rect 273260 3256 273312 3262
rect 273260 3198 273312 3204
rect 273640 480 273668 9250
rect 274652 3330 274680 97974
rect 275204 97866 275232 102037
rect 274744 97838 275232 97866
rect 274744 6662 274772 97838
rect 275756 84194 275784 102037
rect 276216 98002 276244 102037
rect 274836 84166 275784 84194
rect 276032 97974 276244 98002
rect 274836 13258 274864 84166
rect 274824 13252 274876 13258
rect 274824 13194 274876 13200
rect 276032 6914 276060 97974
rect 276676 97866 276704 102037
rect 276124 97838 276704 97866
rect 276124 8906 276152 97838
rect 277136 84194 277164 102037
rect 277688 97968 277716 102037
rect 276216 84166 277164 84194
rect 277412 97940 277716 97968
rect 276216 13190 276244 84166
rect 276204 13184 276256 13190
rect 276204 13126 276256 13132
rect 277124 9240 277176 9246
rect 277124 9182 277176 9188
rect 276112 8900 276164 8906
rect 276112 8842 276164 8848
rect 276032 6886 276152 6914
rect 274732 6656 274784 6662
rect 274732 6598 274784 6604
rect 274824 3936 274876 3942
rect 274824 3878 274876 3884
rect 274640 3324 274692 3330
rect 274640 3266 274692 3272
rect 274836 480 274864 3878
rect 276020 3596 276072 3602
rect 276020 3538 276072 3544
rect 276032 480 276060 3538
rect 276124 3398 276152 6886
rect 276112 3392 276164 3398
rect 276112 3334 276164 3340
rect 277136 480 277164 9182
rect 277412 4146 277440 97940
rect 278148 97866 278176 102037
rect 277504 97838 278176 97866
rect 277504 6594 277532 97838
rect 278608 84194 278636 102037
rect 279160 97968 279188 102037
rect 277596 84166 278636 84194
rect 278792 97940 279188 97968
rect 277596 13122 277624 84166
rect 277584 13116 277636 13122
rect 277584 13058 277636 13064
rect 277492 6588 277544 6594
rect 277492 6530 277544 6536
rect 277400 4140 277452 4146
rect 277400 4082 277452 4088
rect 278792 4078 278820 97940
rect 279620 97866 279648 102037
rect 278884 97838 279648 97866
rect 278884 9654 278912 97838
rect 280080 84194 280108 102037
rect 280632 97968 280660 102037
rect 278976 84166 280108 84194
rect 280172 97940 280660 97968
rect 278976 20330 279004 84166
rect 278964 20324 279016 20330
rect 278964 20266 279016 20272
rect 278872 9648 278924 9654
rect 278872 9590 278924 9596
rect 278780 4072 278832 4078
rect 278780 4014 278832 4020
rect 280172 4010 280200 97940
rect 281092 84194 281120 102037
rect 281552 97968 281580 102037
rect 281552 97940 281764 97968
rect 281632 97844 281684 97850
rect 281632 97786 281684 97792
rect 281540 97776 281592 97782
rect 281540 97718 281592 97724
rect 280264 84166 281120 84194
rect 280264 9586 280292 84166
rect 280252 9580 280304 9586
rect 280252 9522 280304 9528
rect 280712 9172 280764 9178
rect 280712 9114 280764 9120
rect 280160 4004 280212 4010
rect 280160 3946 280212 3952
rect 278320 3868 278372 3874
rect 278320 3810 278372 3816
rect 278332 480 278360 3810
rect 279516 3664 279568 3670
rect 279516 3606 279568 3612
rect 279528 480 279556 3606
rect 280724 480 280752 9114
rect 281552 3942 281580 97718
rect 281644 9518 281672 97786
rect 281736 20262 281764 97940
rect 282012 97782 282040 102037
rect 282564 97850 282592 102037
rect 282920 97980 282972 97986
rect 283024 97968 283052 102037
rect 283484 97986 283512 102037
rect 283472 97980 283524 97986
rect 283024 97940 283144 97968
rect 282920 97922 282972 97928
rect 282552 97844 282604 97850
rect 282552 97786 282604 97792
rect 282000 97776 282052 97782
rect 282000 97718 282052 97724
rect 281724 20256 281776 20262
rect 281724 20198 281776 20204
rect 281632 9512 281684 9518
rect 281632 9454 281684 9460
rect 281540 3936 281592 3942
rect 281540 3878 281592 3884
rect 282932 3874 282960 97922
rect 283012 97844 283064 97850
rect 283012 97786 283064 97792
rect 283024 9450 283052 97786
rect 283116 20194 283144 97940
rect 283472 97922 283524 97928
rect 284036 97850 284064 102037
rect 284392 98048 284444 98054
rect 284392 97990 284444 97996
rect 284300 97980 284352 97986
rect 284300 97922 284352 97928
rect 284024 97844 284076 97850
rect 284024 97786 284076 97792
rect 283104 20188 283156 20194
rect 283104 20130 283156 20136
rect 284312 11490 284340 97922
rect 284300 11484 284352 11490
rect 284300 11426 284352 11432
rect 283012 9444 283064 9450
rect 283012 9386 283064 9392
rect 284300 9104 284352 9110
rect 284300 9046 284352 9052
rect 283104 5772 283156 5778
rect 283104 5714 283156 5720
rect 282920 3868 282972 3874
rect 282920 3810 282972 3816
rect 281908 3800 281960 3806
rect 281908 3742 281960 3748
rect 281920 480 281948 3742
rect 283116 480 283144 5714
rect 284312 480 284340 9046
rect 284404 6526 284432 97990
rect 284496 20126 284524 102037
rect 284956 97986 284984 102037
rect 285416 98054 285444 102037
rect 285772 99680 285824 99686
rect 285772 99622 285824 99628
rect 285404 98048 285456 98054
rect 285404 97990 285456 97996
rect 284944 97980 284996 97986
rect 284944 97922 284996 97928
rect 285680 97980 285732 97986
rect 285680 97922 285732 97928
rect 284484 20120 284536 20126
rect 284484 20062 284536 20068
rect 284484 11484 284536 11490
rect 284484 11426 284536 11432
rect 284392 6520 284444 6526
rect 284392 6462 284444 6468
rect 284496 3806 284524 11426
rect 285404 5296 285456 5302
rect 285404 5238 285456 5244
rect 284484 3800 284536 3806
rect 284484 3742 284536 3748
rect 285416 480 285444 5238
rect 285692 3738 285720 97922
rect 285784 9382 285812 99622
rect 285968 84194 285996 102037
rect 286428 97986 286456 102037
rect 286888 99686 286916 102037
rect 286876 99680 286928 99686
rect 286876 99622 286928 99628
rect 287060 98660 287112 98666
rect 287060 98602 287112 98608
rect 286416 97980 286468 97986
rect 286416 97922 286468 97928
rect 285876 84166 285996 84194
rect 285876 20058 285904 84166
rect 285864 20052 285916 20058
rect 285864 19994 285916 20000
rect 285772 9376 285824 9382
rect 285772 9318 285824 9324
rect 286600 4752 286652 4758
rect 286600 4694 286652 4700
rect 285680 3732 285732 3738
rect 285680 3674 285732 3680
rect 286612 480 286640 4694
rect 287072 3670 287100 98602
rect 287152 97980 287204 97986
rect 287152 97922 287204 97928
rect 287164 9314 287192 97922
rect 287440 84194 287468 102037
rect 287900 98666 287928 102037
rect 287888 98660 287940 98666
rect 287888 98602 287940 98608
rect 288360 97986 288388 102037
rect 288440 100428 288492 100434
rect 288440 100370 288492 100376
rect 288348 97980 288400 97986
rect 288348 97922 288400 97928
rect 287256 84166 287468 84194
rect 287256 14346 287284 84166
rect 287244 14340 287296 14346
rect 287244 14282 287296 14288
rect 287152 9308 287204 9314
rect 287152 9250 287204 9256
rect 287796 9036 287848 9042
rect 287796 8978 287848 8984
rect 287060 3664 287112 3670
rect 287060 3606 287112 3612
rect 287808 480 287836 8978
rect 288452 3534 288480 100370
rect 288912 84194 288940 102037
rect 289372 100434 289400 102037
rect 289360 100428 289412 100434
rect 289360 100370 289412 100376
rect 289832 98002 289860 102037
rect 289832 97974 290044 98002
rect 289912 97912 289964 97918
rect 289912 97854 289964 97860
rect 289820 97844 289872 97850
rect 289820 97786 289872 97792
rect 288544 84166 288940 84194
rect 288544 14414 288572 84166
rect 288532 14408 288584 14414
rect 288532 14350 288584 14356
rect 289832 9246 289860 97786
rect 289924 15162 289952 97854
rect 290016 17814 290044 97974
rect 290292 97850 290320 102037
rect 290844 97918 290872 102037
rect 291304 98002 291332 102037
rect 291200 97980 291252 97986
rect 291304 97974 291424 98002
rect 291764 97986 291792 102037
rect 291200 97922 291252 97928
rect 290832 97912 290884 97918
rect 290832 97854 290884 97860
rect 290280 97844 290332 97850
rect 290280 97786 290332 97792
rect 290004 17808 290056 17814
rect 290004 17750 290056 17756
rect 289912 15156 289964 15162
rect 289912 15098 289964 15104
rect 289820 9240 289872 9246
rect 289820 9182 289872 9188
rect 291212 9178 291240 97922
rect 291292 97912 291344 97918
rect 291292 97854 291344 97860
rect 291304 15094 291332 97854
rect 291396 17746 291424 97974
rect 291752 97980 291804 97986
rect 291752 97922 291804 97928
rect 292316 97918 292344 102037
rect 292672 98048 292724 98054
rect 292672 97990 292724 97996
rect 292580 97980 292632 97986
rect 292580 97922 292632 97928
rect 292304 97912 292356 97918
rect 292304 97854 292356 97860
rect 291384 17740 291436 17746
rect 291384 17682 291436 17688
rect 291292 15088 291344 15094
rect 291292 15030 291344 15036
rect 291200 9172 291252 9178
rect 291200 9114 291252 9120
rect 292592 9110 292620 97922
rect 292684 15026 292712 97990
rect 292776 17678 292804 102037
rect 293236 97986 293264 102037
rect 293696 98054 293724 102037
rect 293684 98048 293736 98054
rect 293684 97990 293736 97996
rect 294052 98048 294104 98054
rect 294052 97990 294104 97996
rect 293224 97980 293276 97986
rect 293224 97922 293276 97928
rect 293960 97980 294012 97986
rect 293960 97922 294012 97928
rect 292764 17672 292816 17678
rect 292764 17614 292816 17620
rect 292672 15020 292724 15026
rect 292672 14962 292724 14968
rect 292580 9104 292632 9110
rect 292580 9046 292632 9052
rect 293972 9042 294000 97922
rect 294064 14958 294092 97990
rect 294248 84194 294276 102037
rect 294708 97986 294736 102037
rect 295168 98054 295196 102037
rect 295156 98048 295208 98054
rect 295156 97990 295208 97996
rect 295432 98048 295484 98054
rect 295432 97990 295484 97996
rect 294696 97980 294748 97986
rect 294696 97922 294748 97928
rect 295340 97980 295392 97986
rect 295340 97922 295392 97928
rect 294156 84166 294276 84194
rect 294156 17610 294184 84166
rect 294144 17604 294196 17610
rect 294144 17546 294196 17552
rect 294052 14952 294104 14958
rect 294052 14894 294104 14900
rect 293960 9036 294012 9042
rect 293960 8978 294012 8984
rect 291384 8968 291436 8974
rect 295352 8945 295380 97922
rect 295444 14822 295472 97990
rect 295720 84194 295748 102037
rect 296180 97986 296208 102037
rect 296640 98054 296668 102037
rect 296628 98048 296680 98054
rect 297100 98002 297128 102037
rect 296628 97990 296680 97996
rect 296168 97980 296220 97986
rect 296168 97922 296220 97928
rect 296732 97974 297128 98002
rect 295536 84166 295748 84194
rect 295536 17542 295564 84166
rect 295524 17536 295576 17542
rect 295524 17478 295576 17484
rect 295432 14816 295484 14822
rect 295432 14758 295484 14764
rect 291384 8910 291436 8916
rect 295338 8936 295394 8945
rect 290188 5500 290240 5506
rect 290188 5442 290240 5448
rect 288992 5228 289044 5234
rect 288992 5170 289044 5176
rect 288440 3528 288492 3534
rect 288440 3470 288492 3476
rect 289004 480 289032 5170
rect 290200 480 290228 5442
rect 291396 480 291424 8910
rect 295338 8871 295394 8880
rect 294880 8628 294932 8634
rect 294880 8570 294932 8576
rect 293684 5840 293736 5846
rect 293684 5782 293736 5788
rect 292580 5092 292632 5098
rect 292580 5034 292632 5040
rect 292592 480 292620 5034
rect 293696 480 293724 5782
rect 294892 480 294920 8570
rect 296076 5160 296128 5166
rect 296076 5102 296128 5108
rect 296088 480 296116 5102
rect 296732 4690 296760 97974
rect 297652 84194 297680 102037
rect 298112 98002 298140 102037
rect 298112 97974 298232 98002
rect 298100 97912 298152 97918
rect 298100 97854 298152 97860
rect 296824 84166 297680 84194
rect 296824 8974 296852 84166
rect 296812 8968 296864 8974
rect 296812 8910 296864 8916
rect 297272 8696 297324 8702
rect 297272 8638 297324 8644
rect 296720 4684 296772 4690
rect 296720 4626 296772 4632
rect 297284 480 297312 8638
rect 298112 4758 298140 97854
rect 298204 14890 298232 97974
rect 298572 97918 298600 102037
rect 298560 97912 298612 97918
rect 298560 97854 298612 97860
rect 299124 84194 299152 102037
rect 299480 97980 299532 97986
rect 299480 97922 299532 97928
rect 298296 84166 299152 84194
rect 298296 19038 298324 84166
rect 298284 19032 298336 19038
rect 298284 18974 298336 18980
rect 298192 14884 298244 14890
rect 298192 14826 298244 14832
rect 298192 10940 298244 10946
rect 298192 10882 298244 10888
rect 298100 4752 298152 4758
rect 298100 4694 298152 4700
rect 203444 354 203472 462
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298204 354 298232 10882
rect 299492 5506 299520 97922
rect 299584 14754 299612 102037
rect 300044 97986 300072 102037
rect 300032 97980 300084 97986
rect 300032 97922 300084 97928
rect 300596 84194 300624 102037
rect 301056 98002 301084 102037
rect 300860 97980 300912 97986
rect 300860 97922 300912 97928
rect 300964 97974 301084 98002
rect 301516 97986 301544 102037
rect 301504 97980 301556 97986
rect 299676 84166 300624 84194
rect 299676 18970 299704 84166
rect 299664 18964 299716 18970
rect 299664 18906 299716 18912
rect 299572 14748 299624 14754
rect 299572 14690 299624 14696
rect 300768 8764 300820 8770
rect 300768 8706 300820 8712
rect 299480 5500 299532 5506
rect 299480 5442 299532 5448
rect 299664 5024 299716 5030
rect 299664 4966 299716 4972
rect 299676 480 299704 4966
rect 300780 480 300808 8706
rect 300872 5438 300900 97922
rect 300964 14686 300992 97974
rect 301504 97922 301556 97928
rect 301976 84194 302004 102037
rect 302528 98002 302556 102037
rect 302240 97980 302292 97986
rect 302240 97922 302292 97928
rect 302344 97974 302556 98002
rect 302988 97986 303016 102037
rect 302976 97980 303028 97986
rect 301056 84166 302004 84194
rect 301056 18902 301084 84166
rect 301044 18896 301096 18902
rect 301044 18838 301096 18844
rect 300952 14680 301004 14686
rect 300952 14622 301004 14628
rect 301504 10872 301556 10878
rect 301504 10814 301556 10820
rect 300860 5432 300912 5438
rect 300860 5374 300912 5380
rect 298438 354 298550 480
rect 298204 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 10814
rect 302252 5370 302280 97922
rect 302344 14618 302372 97974
rect 302976 97922 303028 97928
rect 303448 84194 303476 102037
rect 304000 98002 304028 102037
rect 303620 97980 303672 97986
rect 303620 97922 303672 97928
rect 303724 97974 304028 98002
rect 304460 97986 304488 102037
rect 304448 97980 304500 97986
rect 302436 84166 303476 84194
rect 302436 18834 302464 84166
rect 302424 18828 302476 18834
rect 302424 18770 302476 18776
rect 302332 14612 302384 14618
rect 302332 14554 302384 14560
rect 302240 5364 302292 5370
rect 302240 5306 302292 5312
rect 303632 5302 303660 97922
rect 303724 14550 303752 97974
rect 304448 97922 304500 97928
rect 304920 84194 304948 102037
rect 305000 99952 305052 99958
rect 305000 99894 305052 99900
rect 303816 84166 304948 84194
rect 303816 18766 303844 84166
rect 303804 18760 303856 18766
rect 303804 18702 303856 18708
rect 303896 15904 303948 15910
rect 303896 15846 303948 15852
rect 303712 14544 303764 14550
rect 303712 14486 303764 14492
rect 303620 5296 303672 5302
rect 303620 5238 303672 5244
rect 303160 4956 303212 4962
rect 303160 4898 303212 4904
rect 303172 480 303200 4898
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 15846
rect 305012 5234 305040 99894
rect 305380 84194 305408 102037
rect 305932 99958 305960 102037
rect 305920 99952 305972 99958
rect 305920 99894 305972 99900
rect 306392 98002 306420 102037
rect 306392 97974 306512 98002
rect 306380 97912 306432 97918
rect 306380 97854 306432 97860
rect 305104 84166 305408 84194
rect 305104 14482 305132 84166
rect 305092 14476 305144 14482
rect 305092 14418 305144 14424
rect 305552 10804 305604 10810
rect 305552 10746 305604 10752
rect 305000 5228 305052 5234
rect 305000 5170 305052 5176
rect 305564 480 305592 10746
rect 306392 5166 306420 97854
rect 306484 10198 306512 97974
rect 306852 84194 306880 102037
rect 307404 97918 307432 102037
rect 307760 97980 307812 97986
rect 307760 97922 307812 97928
rect 307392 97912 307444 97918
rect 307392 97854 307444 97860
rect 306576 84166 306880 84194
rect 306576 14521 306604 84166
rect 306562 14512 306618 14521
rect 306562 14447 306618 14456
rect 306472 10192 306524 10198
rect 306472 10134 306524 10140
rect 306380 5160 306432 5166
rect 306380 5102 306432 5108
rect 307772 5098 307800 97922
rect 307864 10266 307892 102037
rect 308324 84194 308352 102037
rect 308784 97986 308812 102037
rect 309336 98002 309364 102037
rect 308772 97980 308824 97986
rect 308772 97922 308824 97928
rect 309140 97980 309192 97986
rect 309140 97922 309192 97928
rect 309244 97974 309364 98002
rect 307956 84166 308352 84194
rect 307956 19990 307984 84166
rect 307944 19984 307996 19990
rect 307944 19926 307996 19932
rect 307944 10736 307996 10742
rect 307944 10678 307996 10684
rect 307852 10260 307904 10266
rect 307852 10202 307904 10208
rect 307760 5092 307812 5098
rect 307760 5034 307812 5040
rect 306748 4888 306800 4894
rect 306748 4830 306800 4836
rect 306760 480 306788 4830
rect 307956 480 307984 10678
rect 309048 10668 309100 10674
rect 309048 10610 309100 10616
rect 309060 480 309088 10610
rect 309152 5030 309180 97922
rect 309244 11014 309272 97974
rect 309796 84194 309824 102037
rect 310256 97986 310284 102037
rect 310808 98002 310836 102037
rect 310244 97980 310296 97986
rect 310244 97922 310296 97928
rect 310520 97980 310572 97986
rect 310520 97922 310572 97928
rect 310624 97974 310836 98002
rect 309336 84166 309824 84194
rect 309336 21554 309364 84166
rect 309324 21548 309376 21554
rect 309324 21490 309376 21496
rect 309232 11008 309284 11014
rect 309232 10950 309284 10956
rect 309140 5024 309192 5030
rect 309140 4966 309192 4972
rect 310532 4962 310560 97922
rect 310624 10946 310652 97974
rect 311268 84194 311296 102037
rect 311728 97986 311756 102037
rect 312280 98002 312308 102037
rect 311716 97980 311768 97986
rect 311716 97922 311768 97928
rect 311900 97980 311952 97986
rect 311900 97922 311952 97928
rect 312004 97974 312308 98002
rect 310716 84166 311296 84194
rect 310716 21486 310744 84166
rect 310704 21480 310756 21486
rect 310704 21422 310756 21428
rect 310612 10940 310664 10946
rect 310612 10882 310664 10888
rect 311440 10600 311492 10606
rect 311440 10542 311492 10548
rect 310520 4956 310572 4962
rect 310520 4898 310572 4904
rect 310242 4856 310298 4865
rect 310242 4791 310298 4800
rect 310256 480 310284 4791
rect 311452 480 311480 10542
rect 311912 4865 311940 97922
rect 312004 10878 312032 97974
rect 312740 84194 312768 102037
rect 313200 97986 313228 102037
rect 313660 98002 313688 102037
rect 313188 97980 313240 97986
rect 313188 97922 313240 97928
rect 313292 97974 313688 98002
rect 312096 84166 312768 84194
rect 312096 21418 312124 84166
rect 312084 21412 312136 21418
rect 312084 21354 312136 21360
rect 311992 10872 312044 10878
rect 311992 10814 312044 10820
rect 313292 10810 313320 97974
rect 314212 84194 314240 102037
rect 313384 84166 314240 84194
rect 313384 16522 313412 84166
rect 313372 16516 313424 16522
rect 313372 16458 313424 16464
rect 313280 10804 313332 10810
rect 313280 10746 313332 10752
rect 312176 10532 312228 10538
rect 312176 10474 312228 10480
rect 311898 4856 311954 4865
rect 311898 4791 311954 4800
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 354 312216 10474
rect 314672 4894 314700 102037
rect 315132 98002 315160 102037
rect 314764 97974 315160 98002
rect 314764 10742 314792 97974
rect 315684 84194 315712 102037
rect 316144 98002 316172 102037
rect 314856 84166 315712 84194
rect 316052 97974 316172 98002
rect 314856 16454 314884 84166
rect 314844 16448 314896 16454
rect 314844 16390 314896 16396
rect 314752 10736 314804 10742
rect 314752 10678 314804 10684
rect 314752 10464 314804 10470
rect 314752 10406 314804 10412
rect 314660 4888 314712 4894
rect 314660 4830 314712 4836
rect 313832 4820 313884 4826
rect 313832 4762 313884 4768
rect 313844 480 313872 4762
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314764 354 314792 10406
rect 316052 4826 316080 97974
rect 316604 97866 316632 102037
rect 316144 97838 316632 97866
rect 316144 10674 316172 97838
rect 317064 84194 317092 102037
rect 317512 98048 317564 98054
rect 317512 97990 317564 97996
rect 317420 97980 317472 97986
rect 317420 97922 317472 97928
rect 316236 84166 317092 84194
rect 316236 16386 316264 84166
rect 316224 16380 316276 16386
rect 316224 16322 316276 16328
rect 316132 10668 316184 10674
rect 316132 10610 316184 10616
rect 317432 10606 317460 97922
rect 317524 16318 317552 97990
rect 317616 17474 317644 102037
rect 318076 97986 318104 102037
rect 318536 98054 318564 102037
rect 318524 98048 318576 98054
rect 318524 97990 318576 97996
rect 318892 98048 318944 98054
rect 318892 97990 318944 97996
rect 318064 97980 318116 97986
rect 318064 97922 318116 97928
rect 318800 97980 318852 97986
rect 318800 97922 318852 97928
rect 317604 17468 317656 17474
rect 317604 17410 317656 17416
rect 317512 16312 317564 16318
rect 317512 16254 317564 16260
rect 317420 10600 317472 10606
rect 317420 10542 317472 10548
rect 318812 10538 318840 97922
rect 318904 16250 318932 97990
rect 319088 84194 319116 102037
rect 319548 97986 319576 102037
rect 320008 98054 320036 102037
rect 319996 98048 320048 98054
rect 319996 97990 320048 97996
rect 320272 98048 320324 98054
rect 320272 97990 320324 97996
rect 319536 97980 319588 97986
rect 319536 97922 319588 97928
rect 320180 97980 320232 97986
rect 320180 97922 320232 97928
rect 318996 84166 319116 84194
rect 318996 17406 319024 84166
rect 318984 17400 319036 17406
rect 318984 17342 319036 17348
rect 318892 16244 318944 16250
rect 318892 16186 318944 16192
rect 318800 10532 318852 10538
rect 318800 10474 318852 10480
rect 320192 10470 320220 97922
rect 320284 11665 320312 97990
rect 320468 84194 320496 102037
rect 321020 97986 321048 102037
rect 321480 98054 321508 102037
rect 321468 98048 321520 98054
rect 321468 97990 321520 97996
rect 321008 97980 321060 97986
rect 321008 97922 321060 97928
rect 321560 97980 321612 97986
rect 321560 97922 321612 97928
rect 320376 84166 320496 84194
rect 320376 17338 320404 84166
rect 320364 17332 320416 17338
rect 320364 17274 320416 17280
rect 320270 11656 320326 11665
rect 320270 11591 320326 11600
rect 320180 10464 320232 10470
rect 320180 10406 320232 10412
rect 318064 10396 318116 10402
rect 318064 10338 318116 10344
rect 316224 10328 316276 10334
rect 316224 10270 316276 10276
rect 316040 4820 316092 4826
rect 316040 4762 316092 4768
rect 316236 480 316264 10270
rect 317328 4548 317380 4554
rect 317328 4490 317380 4496
rect 317340 480 317368 4490
rect 314998 354 315110 480
rect 314764 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 10338
rect 321572 10305 321600 97922
rect 321940 84194 321968 102037
rect 322492 97986 322520 102037
rect 322952 98002 322980 102037
rect 322480 97980 322532 97986
rect 322952 97974 323164 98002
rect 322480 97922 322532 97928
rect 323032 97912 323084 97918
rect 323032 97854 323084 97860
rect 322940 97844 322992 97850
rect 322940 97786 322992 97792
rect 321664 84166 321968 84194
rect 321664 17270 321692 84166
rect 321652 17264 321704 17270
rect 321652 17206 321704 17212
rect 321558 10296 321614 10305
rect 321558 10231 321614 10240
rect 319720 9920 319772 9926
rect 319720 9862 319772 9868
rect 319732 480 319760 9862
rect 322952 6458 322980 97786
rect 323044 10402 323072 97854
rect 323136 16182 323164 97974
rect 323412 97850 323440 102037
rect 323964 97918 323992 102037
rect 324424 98002 324452 102037
rect 324320 97980 324372 97986
rect 324424 97974 324544 98002
rect 324884 97986 324912 102037
rect 324320 97922 324372 97928
rect 323952 97912 324004 97918
rect 323952 97854 324004 97860
rect 323400 97844 323452 97850
rect 323400 97786 323452 97792
rect 323124 16176 323176 16182
rect 323124 16118 323176 16124
rect 323032 10396 323084 10402
rect 323032 10338 323084 10344
rect 323032 9988 323084 9994
rect 323032 9930 323084 9936
rect 322940 6452 322992 6458
rect 322940 6394 322992 6400
rect 322112 6248 322164 6254
rect 322112 6190 322164 6196
rect 320916 4616 320968 4622
rect 320916 4558 320968 4564
rect 320928 480 320956 4558
rect 322124 480 322152 6190
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323044 354 323072 9930
rect 324332 6390 324360 97922
rect 324412 97912 324464 97918
rect 324412 97854 324464 97860
rect 324424 10334 324452 97854
rect 324516 16114 324544 97974
rect 324872 97980 324924 97986
rect 324872 97922 324924 97928
rect 325344 97918 325372 102037
rect 325700 100836 325752 100842
rect 325700 100778 325752 100784
rect 325332 97912 325384 97918
rect 325332 97854 325384 97860
rect 324504 16108 324556 16114
rect 324504 16050 324556 16056
rect 324412 10328 324464 10334
rect 324412 10270 324464 10276
rect 324412 10056 324464 10062
rect 324412 9998 324464 10004
rect 324320 6384 324372 6390
rect 324320 6326 324372 6332
rect 324320 6180 324372 6186
rect 324320 6122 324372 6128
rect 324332 3074 324360 6122
rect 324424 3466 324452 9998
rect 325712 6322 325740 100778
rect 325896 98002 325924 102037
rect 326356 100842 326384 102037
rect 326344 100836 326396 100842
rect 326344 100778 326396 100784
rect 325804 97974 325924 98002
rect 325804 16046 325832 97974
rect 326816 84194 326844 102037
rect 327368 98002 327396 102037
rect 327080 97980 327132 97986
rect 327080 97922 327132 97928
rect 327184 97974 327396 98002
rect 327828 97986 327856 102037
rect 327816 97980 327868 97986
rect 325896 84166 326844 84194
rect 325896 18698 325924 84166
rect 325884 18692 325936 18698
rect 325884 18634 325936 18640
rect 325792 16040 325844 16046
rect 325792 15982 325844 15988
rect 326344 11552 326396 11558
rect 326344 11494 326396 11500
rect 325700 6316 325752 6322
rect 325700 6258 325752 6264
rect 324412 3460 324464 3466
rect 324412 3402 324464 3408
rect 325608 3460 325660 3466
rect 325608 3402 325660 3408
rect 324332 3046 324452 3074
rect 324424 480 324452 3046
rect 325620 480 325648 3402
rect 323278 354 323390 480
rect 323044 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 11494
rect 327092 6254 327120 97922
rect 327184 15978 327212 97974
rect 327816 97922 327868 97928
rect 328288 84194 328316 102037
rect 328748 98002 328776 102037
rect 328460 97980 328512 97986
rect 328460 97922 328512 97928
rect 328564 97974 328776 98002
rect 329300 97986 329328 102037
rect 329288 97980 329340 97986
rect 327276 84166 328316 84194
rect 327276 18630 327304 84166
rect 327264 18624 327316 18630
rect 327264 18566 327316 18572
rect 327172 15972 327224 15978
rect 327172 15914 327224 15920
rect 327080 6248 327132 6254
rect 327080 6190 327132 6196
rect 328472 6186 328500 97922
rect 328564 15910 328592 97974
rect 329288 97922 329340 97928
rect 329760 84194 329788 102037
rect 329840 100972 329892 100978
rect 329840 100914 329892 100920
rect 328656 84166 329788 84194
rect 328656 18601 328684 84166
rect 328642 18592 328698 18601
rect 328642 18527 328698 18536
rect 328552 15904 328604 15910
rect 328552 15846 328604 15852
rect 328736 10124 328788 10130
rect 328736 10066 328788 10072
rect 328460 6180 328512 6186
rect 328460 6122 328512 6128
rect 328000 5908 328052 5914
rect 328000 5850 328052 5856
rect 328012 480 328040 5850
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 10066
rect 329852 3194 329880 100914
rect 330220 84194 330248 102037
rect 330772 100978 330800 102037
rect 330760 100972 330812 100978
rect 330760 100914 330812 100920
rect 329944 84166 330248 84194
rect 329944 15881 329972 84166
rect 329930 15872 329986 15881
rect 329930 15807 329986 15816
rect 330392 14272 330444 14278
rect 330392 14214 330444 14220
rect 329840 3188 329892 3194
rect 329840 3130 329892 3136
rect 330404 480 330432 14214
rect 331232 3602 331260 102037
rect 331692 100434 331720 102068
rect 333244 100496 333296 100502
rect 333244 100438 333296 100444
rect 331680 100428 331732 100434
rect 331680 100370 331732 100376
rect 332600 18420 332652 18426
rect 332600 18362 332652 18368
rect 331588 5976 331640 5982
rect 331588 5918 331640 5924
rect 331220 3596 331272 3602
rect 331220 3538 331272 3544
rect 331600 480 331628 5918
rect 332612 3346 332640 18362
rect 332692 15700 332744 15706
rect 332692 15642 332744 15648
rect 332704 3466 332732 15642
rect 333256 5982 333284 100438
rect 406384 100428 406436 100434
rect 406384 100370 406436 100376
rect 390560 100360 390612 100366
rect 390560 100302 390612 100308
rect 361580 22092 361632 22098
rect 361580 22034 361632 22040
rect 357440 21344 357492 21350
rect 357440 21286 357492 21292
rect 354680 21276 354732 21282
rect 354680 21218 354732 21224
rect 350540 21208 350592 21214
rect 350540 21150 350592 21156
rect 347780 19848 347832 19854
rect 347780 19790 347832 19796
rect 339500 19780 339552 19786
rect 339500 19722 339552 19728
rect 335360 18488 335412 18494
rect 335360 18430 335412 18436
rect 335372 16574 335400 18430
rect 335372 16546 336320 16574
rect 335084 6044 335136 6050
rect 335084 5986 335136 5992
rect 333244 5976 333296 5982
rect 333244 5918 333296 5924
rect 332692 3460 332744 3466
rect 332692 3402 332744 3408
rect 333888 3460 333940 3466
rect 333888 3402 333940 3408
rect 333980 3460 334032 3466
rect 333980 3402 334032 3408
rect 332612 3318 332732 3346
rect 332704 480 332732 3318
rect 333900 480 333928 3402
rect 333992 3194 334020 3402
rect 333980 3188 334032 3194
rect 333980 3130 334032 3136
rect 335096 480 335124 5986
rect 336292 480 336320 16546
rect 337016 15768 337068 15774
rect 337016 15710 337068 15716
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337028 354 337056 15710
rect 338672 6112 338724 6118
rect 338672 6054 338724 6060
rect 338684 480 338712 6054
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 19722
rect 344560 16584 344612 16590
rect 347792 16574 347820 19790
rect 350552 16574 350580 21150
rect 354692 16574 354720 21218
rect 356060 17060 356112 17066
rect 356060 17002 356112 17008
rect 356072 16574 356100 17002
rect 347792 16546 348096 16574
rect 350552 16546 351224 16574
rect 354692 16546 355272 16574
rect 356072 16546 356376 16574
rect 344560 16526 344612 16532
rect 340972 15836 341024 15842
rect 340972 15778 341024 15784
rect 340984 480 341012 15778
rect 342904 11620 342956 11626
rect 342904 11562 342956 11568
rect 342168 6860 342220 6866
rect 342168 6802 342220 6808
rect 342180 480 342208 6802
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 11562
rect 344572 480 344600 16526
rect 346952 11688 347004 11694
rect 346952 11630 347004 11636
rect 345756 6792 345808 6798
rect 345756 6734 345808 6740
rect 345768 480 345796 6734
rect 346964 480 346992 11630
rect 348068 480 348096 16546
rect 349160 12436 349212 12442
rect 349160 12378 349212 12384
rect 349172 3194 349200 12378
rect 349252 6724 349304 6730
rect 349252 6666 349304 6672
rect 349160 3188 349212 3194
rect 349160 3130 349212 3136
rect 349264 480 349292 6666
rect 350448 3188 350500 3194
rect 350448 3130 350500 3136
rect 350460 480 350488 3130
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 353576 12368 353628 12374
rect 353576 12310 353628 12316
rect 352838 6216 352894 6225
rect 352838 6151 352894 6160
rect 352852 480 352880 6151
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 12310
rect 355244 480 355272 16546
rect 356348 480 356376 16546
rect 357452 3194 357480 21286
rect 358820 17128 358872 17134
rect 358820 17070 358872 17076
rect 358832 16574 358860 17070
rect 361592 16574 361620 22034
rect 365720 22024 365772 22030
rect 365720 21966 365772 21972
rect 362960 17196 363012 17202
rect 362960 17138 363012 17144
rect 362972 16574 363000 17138
rect 358832 16546 359504 16574
rect 361592 16546 361896 16574
rect 362972 16546 363552 16574
rect 357532 12300 357584 12306
rect 357532 12242 357584 12248
rect 357440 3188 357492 3194
rect 357440 3130 357492 3136
rect 357544 480 357572 12242
rect 358728 3188 358780 3194
rect 358728 3130 358780 3136
rect 358740 480 358768 3130
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 361120 12232 361172 12238
rect 361120 12174 361172 12180
rect 361132 480 361160 12174
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363524 480 363552 16546
rect 364616 12164 364668 12170
rect 364616 12106 364668 12112
rect 364628 480 364656 12106
rect 365732 3074 365760 21966
rect 368480 21956 368532 21962
rect 368480 21898 368532 21904
rect 365812 17944 365864 17950
rect 365812 17886 365864 17892
rect 365824 3194 365852 17886
rect 368492 16574 368520 21898
rect 372620 21888 372672 21894
rect 372620 21830 372672 21836
rect 369860 17876 369912 17882
rect 369860 17818 369912 17824
rect 369872 16574 369900 17818
rect 372632 16574 372660 21830
rect 375380 21820 375432 21826
rect 375380 21762 375432 21768
rect 375392 16574 375420 21762
rect 379520 21752 379572 21758
rect 379520 21694 379572 21700
rect 368492 16546 369440 16574
rect 369872 16546 370176 16574
rect 372632 16546 372936 16574
rect 375392 16546 376064 16574
rect 367744 12096 367796 12102
rect 367744 12038 367796 12044
rect 365812 3188 365864 3194
rect 365812 3130 365864 3136
rect 367008 3188 367060 3194
rect 367008 3130 367060 3136
rect 365732 3046 365852 3074
rect 365824 480 365852 3046
rect 367020 480 367048 3130
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 12038
rect 369412 480 369440 16546
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 16546
rect 371240 12028 371292 12034
rect 371240 11970 371292 11976
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 11970
rect 372908 480 372936 16546
rect 374000 11960 374052 11966
rect 374000 11902 374052 11908
rect 374012 3194 374040 11902
rect 374092 7404 374144 7410
rect 374092 7346 374144 7352
rect 374000 3188 374052 3194
rect 374000 3130 374052 3136
rect 374104 480 374132 7346
rect 375288 3188 375340 3194
rect 375288 3130 375340 3136
rect 375300 480 375328 3130
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 378416 11892 378468 11898
rect 378416 11834 378468 11840
rect 377680 7472 377732 7478
rect 377680 7414 377732 7420
rect 377692 480 377720 7414
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 11834
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 21694
rect 382280 21684 382332 21690
rect 382280 21626 382332 21632
rect 381176 7540 381228 7546
rect 381176 7482 381228 7488
rect 381188 480 381216 7482
rect 382292 3194 382320 21626
rect 386420 21616 386472 21622
rect 386420 21558 386472 21564
rect 386432 16574 386460 21558
rect 389180 19916 389232 19922
rect 389180 19858 389232 19864
rect 389192 16574 389220 19858
rect 390572 16574 390600 100302
rect 397460 100292 397512 100298
rect 397460 100234 397512 100240
rect 393320 23180 393372 23186
rect 393320 23122 393372 23128
rect 391940 20596 391992 20602
rect 391940 20538 391992 20544
rect 391952 16574 391980 20538
rect 393332 16574 393360 23122
rect 396080 20528 396132 20534
rect 396080 20470 396132 20476
rect 386432 16546 386736 16574
rect 389192 16546 389496 16574
rect 390572 16546 390692 16574
rect 391952 16546 392624 16574
rect 393332 16546 394280 16574
rect 382372 11824 382424 11830
rect 382372 11766 382424 11772
rect 382280 3188 382332 3194
rect 382280 3130 382332 3136
rect 382384 480 382412 11766
rect 385960 11756 386012 11762
rect 385960 11698 386012 11704
rect 384764 8288 384816 8294
rect 384764 8230 384816 8236
rect 383568 3188 383620 3194
rect 383568 3130 383620 3136
rect 383580 480 383608 3130
rect 384776 480 384804 8230
rect 385972 480 386000 11698
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 388260 8220 388312 8226
rect 388260 8162 388312 8168
rect 388272 480 388300 8162
rect 389468 480 389496 16546
rect 390664 480 390692 16546
rect 391848 8152 391900 8158
rect 391848 8094 391900 8100
rect 391860 480 391888 8094
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387126 -960 387238 326
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394252 480 394280 16546
rect 395344 8084 395396 8090
rect 395344 8026 395396 8032
rect 395356 480 395384 8026
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 20470
rect 397472 16574 397500 100234
rect 404360 100224 404412 100230
rect 404360 100166 404412 100172
rect 400220 23112 400272 23118
rect 400220 23054 400272 23060
rect 398840 20460 398892 20466
rect 398840 20402 398892 20408
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398852 3194 398880 20402
rect 400232 16574 400260 23054
rect 402980 20392 403032 20398
rect 402980 20334 403032 20340
rect 402992 16574 403020 20334
rect 400232 16546 400904 16574
rect 402992 16546 403664 16574
rect 398932 8016 398984 8022
rect 398932 7958 398984 7964
rect 398840 3188 398892 3194
rect 398840 3130 398892 3136
rect 398944 480 398972 7958
rect 400128 3188 400180 3194
rect 400128 3130 400180 3136
rect 400140 480 400168 3130
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402520 7948 402572 7954
rect 402520 7890 402572 7896
rect 402532 480 402560 7890
rect 403636 480 403664 16546
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 100166
rect 406016 7880 406068 7886
rect 406016 7822 406068 7828
rect 406028 480 406056 7822
rect 406396 3369 406424 100370
rect 411260 100156 411312 100162
rect 411260 100098 411312 100104
rect 407120 23044 407172 23050
rect 407120 22986 407172 22992
rect 406382 3360 406438 3369
rect 406382 3295 406438 3304
rect 407132 3194 407160 22986
rect 411272 16574 411300 100098
rect 425060 100088 425112 100094
rect 425060 100030 425112 100036
rect 415400 22976 415452 22982
rect 415400 22918 415452 22924
rect 415412 16574 415440 22918
rect 422300 22908 422352 22914
rect 422300 22850 422352 22856
rect 422312 16574 422340 22850
rect 423680 18556 423732 18562
rect 423680 18498 423732 18504
rect 411272 16546 411944 16574
rect 415412 16546 415532 16574
rect 422312 16546 422616 16574
rect 410800 12980 410852 12986
rect 410800 12922 410852 12928
rect 407212 12912 407264 12918
rect 407212 12854 407264 12860
rect 407120 3188 407172 3194
rect 407120 3130 407172 3136
rect 407224 480 407252 12854
rect 409604 7812 409656 7818
rect 409604 7754 409656 7760
rect 408408 3188 408460 3194
rect 408408 3130 408460 3136
rect 408420 480 408448 3130
rect 409616 480 409644 7754
rect 410812 480 410840 12922
rect 411916 480 411944 16546
rect 414296 13048 414348 13054
rect 414296 12990 414348 12996
rect 413100 7744 413152 7750
rect 413100 7686 413152 7692
rect 413112 480 413140 7686
rect 414308 480 414336 12990
rect 415504 480 415532 16546
rect 417424 13796 417476 13802
rect 417424 13738 417476 13744
rect 416688 7676 416740 7682
rect 416688 7618 416740 7624
rect 416700 480 416728 7618
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 13738
rect 420920 13728 420972 13734
rect 420920 13670 420972 13676
rect 420184 7608 420236 7614
rect 420184 7550 420236 7556
rect 418988 5976 419040 5982
rect 418988 5918 419040 5924
rect 419000 480 419028 5918
rect 420196 480 420224 7550
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 417854 -960 417966 326
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 354 420960 13670
rect 422588 480 422616 16546
rect 423692 3074 423720 18498
rect 425072 16574 425100 100030
rect 431960 100020 432012 100026
rect 431960 99962 432012 99968
rect 429200 22840 429252 22846
rect 429200 22782 429252 22788
rect 426440 19304 426492 19310
rect 426440 19246 426492 19252
rect 426452 16574 426480 19246
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 423772 13660 423824 13666
rect 423772 13602 423824 13608
rect 423784 3194 423812 13602
rect 423772 3188 423824 3194
rect 423772 3130 423824 3136
rect 424968 3188 425020 3194
rect 424968 3130 425020 3136
rect 423692 3046 423812 3074
rect 423784 480 423812 3046
rect 424980 480 425008 3130
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428464 13592 428516 13598
rect 428464 13534 428516 13540
rect 428476 480 428504 13534
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 22782
rect 430580 19236 430632 19242
rect 430580 19178 430632 19184
rect 430592 16574 430620 19178
rect 430592 16546 430896 16574
rect 430868 480 430896 16546
rect 431972 3194 432000 99962
rect 577516 33114 577544 343674
rect 577608 73166 577636 343742
rect 577700 100706 577728 347754
rect 580264 343868 580316 343874
rect 580264 343810 580316 343816
rect 579618 343768 579674 343777
rect 579618 343703 579674 343712
rect 579632 343670 579660 343703
rect 579620 343664 579672 343670
rect 579620 343606 579672 343612
rect 580080 341080 580132 341086
rect 580080 341022 580132 341028
rect 580092 325281 580120 341022
rect 580172 340944 580224 340950
rect 580172 340886 580224 340892
rect 580078 325272 580134 325281
rect 580078 325207 580134 325216
rect 580080 272604 580132 272610
rect 580080 272546 580132 272552
rect 580092 232393 580120 272546
rect 580184 245585 580212 340886
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580078 232384 580134 232393
rect 580078 232319 580134 232328
rect 577688 100700 577740 100706
rect 577688 100642 577740 100648
rect 579988 100700 580040 100706
rect 579988 100642 580040 100648
rect 580000 99521 580028 100642
rect 579986 99512 580042 99521
rect 579986 99447 580042 99456
rect 580276 86193 580304 343810
rect 580816 342508 580868 342514
rect 580816 342450 580868 342456
rect 580632 342440 580684 342446
rect 580632 342382 580684 342388
rect 580540 342372 580592 342378
rect 580540 342314 580592 342320
rect 580448 342304 580500 342310
rect 580448 342246 580500 342252
rect 580354 340912 580410 340921
rect 580354 340847 580410 340856
rect 580368 112849 580396 340847
rect 580460 126041 580488 342246
rect 580552 165889 580580 342314
rect 580644 179217 580672 342382
rect 580722 341048 580778 341057
rect 580722 340983 580778 340992
rect 580736 192545 580764 340983
rect 580828 205737 580856 342450
rect 580908 341012 580960 341018
rect 580908 340954 580960 340960
rect 580920 298761 580948 340954
rect 580906 298752 580962 298761
rect 580906 298687 580962 298696
rect 580908 272536 580960 272542
rect 580908 272478 580960 272484
rect 580814 205728 580870 205737
rect 580814 205663 580870 205672
rect 580722 192536 580778 192545
rect 580722 192471 580778 192480
rect 580630 179208 580686 179217
rect 580630 179143 580686 179152
rect 580538 165880 580594 165889
rect 580538 165815 580594 165824
rect 580920 152697 580948 272478
rect 580906 152688 580962 152697
rect 580906 152623 580962 152632
rect 580446 126032 580502 126041
rect 580446 125967 580502 125976
rect 580354 112840 580410 112849
rect 580354 112775 580410 112784
rect 580262 86184 580318 86193
rect 580262 86119 580318 86128
rect 577596 73160 577648 73166
rect 577596 73102 577648 73108
rect 579712 73160 579764 73166
rect 579712 73102 579764 73108
rect 579724 73001 579752 73102
rect 579710 72992 579766 73001
rect 579710 72927 579766 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 579618 33144 579674 33153
rect 577504 33108 577556 33114
rect 579618 33079 579620 33088
rect 577504 33050 577556 33056
rect 579672 33079 579674 33088
rect 579620 33050 579672 33056
rect 436100 22772 436152 22778
rect 436100 22714 436152 22720
rect 433340 19168 433392 19174
rect 433340 19110 433392 19116
rect 433352 16574 433380 19110
rect 436112 16574 436140 22714
rect 528560 21548 528612 21554
rect 528560 21490 528612 21496
rect 456892 20324 456944 20330
rect 456892 20266 456944 20272
rect 437480 19100 437532 19106
rect 437480 19042 437532 19048
rect 433352 16546 434024 16574
rect 436112 16546 436784 16574
rect 432052 13524 432104 13530
rect 432052 13466 432104 13472
rect 431960 3188 432012 3194
rect 431960 3130 432012 3136
rect 432064 480 432092 13466
rect 433248 3188 433300 3194
rect 433248 3130 433300 3136
rect 433260 480 433288 3130
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 435088 13456 435140 13462
rect 435088 13398 435140 13404
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 13398
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 19042
rect 439136 13388 439188 13394
rect 439136 13330 439188 13336
rect 439148 480 439176 13330
rect 442632 13320 442684 13326
rect 442632 13262 442684 13268
rect 441528 8832 441580 8838
rect 441528 8774 441580 8780
rect 440332 3256 440384 3262
rect 440332 3198 440384 3204
rect 440344 480 440372 3198
rect 441540 480 441568 8774
rect 442644 480 442672 13262
rect 445760 13252 445812 13258
rect 445760 13194 445812 13200
rect 445024 6656 445076 6662
rect 445024 6598 445076 6604
rect 443828 3324 443880 3330
rect 443828 3266 443880 3272
rect 443840 480 443868 3266
rect 445036 480 445064 6598
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 13194
rect 448520 13184 448572 13190
rect 448520 13126 448572 13132
rect 448532 3398 448560 13126
rect 453304 13116 453356 13122
rect 453304 13058 453356 13064
rect 448612 8900 448664 8906
rect 448612 8842 448664 8848
rect 447416 3392 447468 3398
rect 447416 3334 447468 3340
rect 448520 3392 448572 3398
rect 448520 3334 448572 3340
rect 447428 480 447456 3334
rect 448624 480 448652 8842
rect 452108 6588 452160 6594
rect 452108 6530 452160 6536
rect 450912 4140 450964 4146
rect 450912 4082 450964 4088
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 449820 480 449848 3334
rect 450924 480 450952 4082
rect 452120 480 452148 6530
rect 453316 480 453344 13058
rect 455696 9648 455748 9654
rect 455696 9590 455748 9596
rect 454500 4072 454552 4078
rect 454500 4014 454552 4020
rect 454512 480 454540 4014
rect 455708 480 455736 9590
rect 456904 480 456932 20266
rect 459560 20256 459612 20262
rect 459560 20198 459612 20204
rect 459572 16574 459600 20198
rect 463700 20188 463752 20194
rect 463700 20130 463752 20136
rect 463712 16574 463740 20130
rect 466460 20120 466512 20126
rect 466460 20062 466512 20068
rect 466472 16574 466500 20062
rect 470600 20052 470652 20058
rect 470600 19994 470652 20000
rect 459572 16546 459968 16574
rect 463712 16546 464016 16574
rect 466472 16546 467512 16574
rect 459192 9580 459244 9586
rect 459192 9522 459244 9528
rect 458088 4004 458140 4010
rect 458088 3946 458140 3952
rect 458100 480 458128 3946
rect 459204 480 459232 9522
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 462780 9512 462832 9518
rect 462780 9454 462832 9460
rect 461584 3936 461636 3942
rect 461584 3878 461636 3884
rect 461596 480 461624 3878
rect 462792 480 462820 9454
rect 463988 480 464016 16546
rect 466276 9444 466328 9450
rect 466276 9386 466328 9392
rect 465172 3868 465224 3874
rect 465172 3810 465224 3816
rect 465184 480 465212 3810
rect 466288 480 466316 9386
rect 467484 480 467512 16546
rect 469864 6520 469916 6526
rect 469864 6462 469916 6468
rect 468668 3800 468720 3806
rect 468668 3742 468720 3748
rect 468680 480 468708 3742
rect 469876 480 469904 6462
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 19994
rect 524420 19984 524472 19990
rect 524420 19926 524472 19932
rect 502340 19032 502392 19038
rect 502340 18974 502392 18980
rect 480260 17808 480312 17814
rect 480260 17750 480312 17756
rect 480272 16574 480300 17750
rect 483020 17740 483072 17746
rect 483020 17682 483072 17688
rect 483032 16574 483060 17682
rect 487160 17672 487212 17678
rect 487160 17614 487212 17620
rect 480272 16546 480576 16574
rect 483032 16546 484072 16574
rect 478144 14408 478196 14414
rect 478144 14350 478196 14356
rect 474096 14340 474148 14346
rect 474096 14282 474148 14288
rect 473452 9376 473504 9382
rect 473452 9318 473504 9324
rect 472256 3732 472308 3738
rect 472256 3674 472308 3680
rect 472268 480 472296 3674
rect 473464 480 473492 9318
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 14282
rect 476948 9308 477000 9314
rect 476948 9250 477000 9256
rect 475752 3664 475804 3670
rect 475752 3606 475804 3612
rect 475764 480 475792 3606
rect 476960 480 476988 9250
rect 478156 480 478184 14350
rect 479340 3528 479392 3534
rect 479340 3470 479392 3476
rect 479352 480 479380 3470
rect 480548 480 480576 16546
rect 482376 15156 482428 15162
rect 482376 15098 482428 15104
rect 481732 9240 481784 9246
rect 481732 9182 481784 9188
rect 481744 480 481772 9182
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 15098
rect 484044 480 484072 16546
rect 486424 15088 486476 15094
rect 486424 15030 486476 15036
rect 485228 9172 485280 9178
rect 485228 9114 485280 9120
rect 485240 480 485268 9114
rect 486436 480 486464 15030
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487172 354 487200 17614
rect 489920 17604 489972 17610
rect 489920 17546 489972 17552
rect 488816 9104 488868 9110
rect 488816 9046 488868 9052
rect 488828 480 488856 9046
rect 489932 3534 489960 17546
rect 494060 17536 494112 17542
rect 494060 17478 494112 17484
rect 494072 16574 494100 17478
rect 502352 16574 502380 18974
rect 506480 18964 506532 18970
rect 506480 18906 506532 18912
rect 494072 16546 494744 16574
rect 502352 16546 503024 16574
rect 490012 15020 490064 15026
rect 490012 14962 490064 14968
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 490024 3346 490052 14962
rect 493048 14952 493100 14958
rect 493048 14894 493100 14900
rect 492312 9036 492364 9042
rect 492312 8978 492364 8984
rect 490748 3528 490800 3534
rect 490748 3470 490800 3476
rect 489932 3318 490052 3346
rect 489932 480 489960 3318
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3470
rect 492324 480 492352 8978
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 14894
rect 494716 480 494744 16546
rect 500592 14884 500644 14890
rect 500592 14826 500644 14832
rect 497096 14816 497148 14822
rect 497096 14758 497148 14764
rect 495898 8936 495954 8945
rect 495898 8871 495954 8880
rect 495912 480 495940 8871
rect 497108 480 497136 14758
rect 499396 8968 499448 8974
rect 499396 8910 499448 8916
rect 498200 4684 498252 4690
rect 498200 4626 498252 4632
rect 498212 480 498240 4626
rect 499408 480 499436 8910
rect 500604 480 500632 14826
rect 501788 4752 501840 4758
rect 501788 4694 501840 4700
rect 501800 480 501828 4694
rect 502996 480 503024 16546
rect 503720 14748 503772 14754
rect 503720 14690 503772 14696
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 14690
rect 505376 5500 505428 5506
rect 505376 5442 505428 5448
rect 505388 480 505416 5442
rect 506492 480 506520 18906
rect 509240 18896 509292 18902
rect 509240 18838 509292 18844
rect 509252 16574 509280 18838
rect 513380 18828 513432 18834
rect 513380 18770 513432 18776
rect 509252 16546 509648 16574
rect 507216 14680 507268 14686
rect 507216 14622 507268 14628
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 14622
rect 508872 5432 508924 5438
rect 508872 5374 508924 5380
rect 508884 480 508912 5374
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511264 14612 511316 14618
rect 511264 14554 511316 14560
rect 511276 480 511304 14554
rect 512460 5364 512512 5370
rect 512460 5306 512512 5312
rect 512472 480 512500 5306
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513392 354 513420 18770
rect 516140 18760 516192 18766
rect 516140 18702 516192 18708
rect 516152 16574 516180 18702
rect 524432 16574 524460 19926
rect 516152 16546 517192 16574
rect 524432 16546 525472 16574
rect 514760 14544 514812 14550
rect 514760 14486 514812 14492
rect 514772 480 514800 14486
rect 515956 5296 516008 5302
rect 515956 5238 516008 5244
rect 515968 480 515996 5238
rect 517164 480 517192 16546
rect 521658 14512 521714 14521
rect 517888 14476 517940 14482
rect 521658 14447 521714 14456
rect 517888 14418 517940 14424
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 14418
rect 520280 10192 520332 10198
rect 520280 10134 520332 10140
rect 519544 5228 519596 5234
rect 519544 5170 519596 5176
rect 519556 480 519584 5170
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 10134
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 14447
rect 523776 10260 523828 10266
rect 523776 10202 523828 10208
rect 523040 5160 523092 5166
rect 523040 5102 523092 5108
rect 523052 480 523080 5102
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 10202
rect 525444 480 525472 16546
rect 527824 11008 527876 11014
rect 527824 10950 527876 10956
rect 526628 5092 526680 5098
rect 526628 5034 526680 5040
rect 526640 480 526668 5034
rect 527836 480 527864 10950
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 354 528600 21490
rect 531320 21480 531372 21486
rect 531320 21422 531372 21428
rect 530124 5024 530176 5030
rect 530124 4966 530176 4972
rect 530136 480 530164 4966
rect 531332 3534 531360 21422
rect 535460 21412 535512 21418
rect 535460 21354 535512 21360
rect 535472 16574 535500 21354
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 569960 18692 570012 18698
rect 569960 18634 570012 18640
rect 547880 17468 547932 17474
rect 547880 17410 547932 17416
rect 535472 16546 536144 16574
rect 531412 10940 531464 10946
rect 531412 10882 531464 10888
rect 531320 3528 531372 3534
rect 531320 3470 531372 3476
rect 531424 3346 531452 10882
rect 534448 10872 534500 10878
rect 534448 10814 534500 10820
rect 533712 4956 533764 4962
rect 533712 4898 533764 4904
rect 532148 3528 532200 3534
rect 532148 3470 532200 3476
rect 531332 3318 531452 3346
rect 531332 480 531360 3318
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 528990 -960 529102 326
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532160 354 532188 3470
rect 533724 480 533752 4898
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 10814
rect 536116 480 536144 16546
rect 539600 16516 539652 16522
rect 539600 16458 539652 16464
rect 538220 10804 538272 10810
rect 538220 10746 538272 10752
rect 537206 4856 537262 4865
rect 537206 4791 537262 4800
rect 537220 480 537248 4791
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 10746
rect 539612 480 539640 16458
rect 542728 16448 542780 16454
rect 542728 16390 542780 16396
rect 541992 10736 542044 10742
rect 541992 10678 542044 10684
rect 540796 4888 540848 4894
rect 540796 4830 540848 4836
rect 540808 480 540836 4830
rect 542004 480 542032 10678
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 354 542768 16390
rect 546500 16380 546552 16386
rect 546500 16322 546552 16328
rect 545488 10668 545540 10674
rect 545488 10610 545540 10616
rect 544384 4820 544436 4826
rect 544384 4762 544436 4768
rect 544396 480 544424 4762
rect 545500 480 545528 10610
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 16322
rect 547892 480 547920 17410
rect 550640 17400 550692 17406
rect 550640 17342 550692 17348
rect 550652 16574 550680 17342
rect 554780 17332 554832 17338
rect 554780 17274 554832 17280
rect 550652 16546 551048 16574
rect 550272 16312 550324 16318
rect 550272 16254 550324 16260
rect 548616 10600 548668 10606
rect 548616 10542 548668 10548
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548628 354 548656 10542
rect 550284 480 550312 16254
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 553768 16244 553820 16250
rect 553768 16186 553820 16192
rect 552664 10532 552716 10538
rect 552664 10474 552716 10480
rect 552676 480 552704 10474
rect 553780 480 553808 16186
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 17274
rect 557540 17264 557592 17270
rect 557540 17206 557592 17212
rect 557552 16574 557580 17206
rect 569972 16574 570000 18634
rect 572720 18624 572772 18630
rect 572720 18566 572772 18572
rect 576858 18592 576914 18601
rect 572732 16574 572760 18566
rect 576858 18527 576914 18536
rect 576872 16574 576900 18527
rect 557552 16546 558592 16574
rect 569972 16546 570368 16574
rect 572732 16546 573496 16574
rect 576872 16546 576992 16574
rect 556158 11656 556214 11665
rect 556158 11591 556214 11600
rect 556172 3534 556200 11591
rect 556252 10464 556304 10470
rect 556252 10406 556304 10412
rect 556160 3528 556212 3534
rect 556160 3470 556212 3476
rect 556264 3346 556292 10406
rect 556988 3528 557040 3534
rect 556988 3470 557040 3476
rect 556172 3318 556292 3346
rect 556172 480 556200 3318
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 557000 354 557028 3470
rect 558564 480 558592 16546
rect 560392 16176 560444 16182
rect 560392 16118 560444 16124
rect 559286 10296 559342 10305
rect 559286 10231 559342 10240
rect 557326 354 557438 480
rect 557000 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 10231
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16118
rect 564440 16108 564492 16114
rect 564440 16050 564492 16056
rect 563060 10396 563112 10402
rect 563060 10338 563112 10344
rect 562048 6452 562100 6458
rect 562048 6394 562100 6400
rect 562060 480 562088 6394
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 10338
rect 564452 480 564480 16050
rect 567568 16040 567620 16046
rect 567568 15982 567620 15988
rect 566832 10328 566884 10334
rect 566832 10270 566884 10276
rect 565636 6384 565688 6390
rect 565636 6326 565688 6332
rect 565648 480 565676 6326
rect 566844 480 566872 10270
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567580 354 567608 15982
rect 569132 6316 569184 6322
rect 569132 6258 569184 6264
rect 569144 480 569172 6258
rect 570340 480 570368 16546
rect 571340 15972 571392 15978
rect 571340 15914 571392 15920
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 15914
rect 572720 6248 572772 6254
rect 572720 6190 572772 6196
rect 572732 480 572760 6190
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 575112 15904 575164 15910
rect 575112 15846 575164 15852
rect 575124 480 575152 15846
rect 576308 6180 576360 6186
rect 576308 6122 576360 6128
rect 576320 480 576348 6122
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 576964 354 576992 16546
rect 578606 15872 578662 15881
rect 578606 15807 578662 15816
rect 578620 480 578648 15807
rect 582196 3596 582248 3602
rect 582196 3538 582248 3544
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 3538
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 671200 3478 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3238 462576 3294 462632
rect 3146 449520 3202 449576
rect 3422 423544 3478 423600
rect 3146 410488 3202 410544
rect 3422 397468 3424 397488
rect 3424 397468 3476 397488
rect 3476 397468 3478 397488
rect 3422 397432 3478 397468
rect 3422 371320 3478 371376
rect 3146 358400 3202 358456
rect 3330 345344 3386 345400
rect 99286 344664 99342 344720
rect 3238 319232 3294 319288
rect 3330 306176 3386 306232
rect 2778 162832 2834 162888
rect 4066 293120 4122 293176
rect 3974 267144 4030 267200
rect 3882 254088 3938 254144
rect 3790 241032 3846 241088
rect 3698 214920 3754 214976
rect 3606 201864 3662 201920
rect 3514 188808 3570 188864
rect 3422 149776 3478 149832
rect 90362 341264 90418 341320
rect 2778 110608 2834 110664
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3146 32408 3202 32464
rect 5262 3304 5318 3360
rect 13542 6160 13598 6216
rect 90546 341400 90602 341456
rect 65522 4800 65578 4856
rect 141422 344528 141478 344584
rect 135074 344392 135130 344448
rect 116122 343984 116178 344040
rect 132958 344256 133014 344312
rect 128818 344120 128874 344176
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 309874 343848 309930 343904
rect 108118 341536 108174 341592
rect 120630 341536 120686 341592
rect 135350 341536 135406 341592
rect 164146 341536 164202 341592
rect 322202 341400 322258 341456
rect 326434 341400 326490 341456
rect 328458 341400 328514 341456
rect 330666 341400 330722 341456
rect 94042 3304 94098 3360
rect 96710 6160 96766 6216
rect 109314 3304 109370 3360
rect 118790 4800 118846 4856
rect 136730 3304 136786 3360
rect 219438 4800 219494 4856
rect 236274 6160 236330 6216
rect 295338 8880 295394 8936
rect 306562 14456 306618 14512
rect 310242 4800 310298 4856
rect 311898 4800 311954 4856
rect 320270 11600 320326 11656
rect 321558 10240 321614 10296
rect 328642 18536 328698 18592
rect 329930 15816 329986 15872
rect 352838 6160 352894 6216
rect 406382 3304 406438 3360
rect 579618 343712 579674 343768
rect 580078 325216 580134 325272
rect 580170 245520 580226 245576
rect 580078 232328 580134 232384
rect 579986 99456 580042 99512
rect 580354 340856 580410 340912
rect 580722 340992 580778 341048
rect 580906 298696 580962 298752
rect 580814 205672 580870 205728
rect 580722 192480 580778 192536
rect 580630 179152 580686 179208
rect 580538 165824 580594 165880
rect 580906 152632 580962 152688
rect 580446 125976 580502 126032
rect 580354 112784 580410 112840
rect 580262 86128 580318 86184
rect 579710 72936 579766 72992
rect 580170 59608 580226 59664
rect 579618 33108 579674 33144
rect 579618 33088 579620 33108
rect 579620 33088 579672 33108
rect 579672 33088 579674 33108
rect 495898 8880 495954 8936
rect 521658 14456 521714 14512
rect 579986 19760 580042 19816
rect 537206 4800 537262 4856
rect 576858 18536 576914 18592
rect 556158 11600 556214 11656
rect 559286 10240 559342 10296
rect 578606 15816 578662 15872
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 99281 344722 99347 344725
rect 580206 344722 580212 344724
rect 99281 344720 580212 344722
rect 99281 344664 99286 344720
rect 99342 344664 580212 344720
rect 99281 344662 580212 344664
rect 99281 344659 99347 344662
rect 580206 344660 580212 344662
rect 580276 344660 580282 344724
rect 141417 344586 141483 344589
rect 328126 344586 328132 344588
rect 141417 344584 328132 344586
rect 141417 344528 141422 344584
rect 141478 344528 328132 344584
rect 141417 344526 328132 344528
rect 141417 344523 141483 344526
rect 328126 344524 328132 344526
rect 328196 344524 328202 344588
rect 135069 344450 135135 344453
rect 327942 344450 327948 344452
rect 135069 344448 327948 344450
rect 135069 344392 135074 344448
rect 135130 344392 327948 344448
rect 135069 344390 327948 344392
rect 135069 344387 135135 344390
rect 327942 344388 327948 344390
rect 328012 344388 328018 344452
rect 132953 344314 133019 344317
rect 329046 344314 329052 344316
rect 132953 344312 329052 344314
rect 132953 344256 132958 344312
rect 133014 344256 329052 344312
rect 132953 344254 329052 344256
rect 132953 344251 133019 344254
rect 329046 344252 329052 344254
rect 329116 344252 329122 344316
rect 128813 344178 128879 344181
rect 327758 344178 327764 344180
rect 128813 344176 327764 344178
rect 128813 344120 128818 344176
rect 128874 344120 327764 344176
rect 128813 344118 327764 344120
rect 128813 344115 128879 344118
rect 327758 344116 327764 344118
rect 327828 344116 327834 344180
rect 116117 344042 116183 344045
rect 327574 344042 327580 344044
rect 116117 344040 327580 344042
rect 116117 343984 116122 344040
rect 116178 343984 327580 344040
rect 116117 343982 327580 343984
rect 116117 343979 116183 343982
rect 327574 343980 327580 343982
rect 327644 343980 327650 344044
rect 3550 343844 3556 343908
rect 3620 343906 3626 343908
rect 309869 343906 309935 343909
rect 3620 343904 309935 343906
rect 3620 343848 309874 343904
rect 309930 343848 309935 343904
rect 3620 343846 309935 343848
rect 3620 343844 3626 343846
rect 309869 343843 309935 343846
rect 579613 343770 579679 343773
rect 580758 343770 580764 343772
rect 579613 343768 580764 343770
rect 579613 343712 579618 343768
rect 579674 343712 580764 343768
rect 579613 343710 580764 343712
rect 579613 343707 579679 343710
rect 580758 343708 580764 343710
rect 580828 343708 580834 343772
rect 108113 341594 108179 341597
rect 110454 341594 110460 341596
rect 108113 341592 110460 341594
rect 108113 341536 108118 341592
rect 108174 341536 110460 341592
rect 108113 341534 110460 341536
rect 108113 341531 108179 341534
rect 110454 341532 110460 341534
rect 110524 341532 110530 341596
rect 120625 341594 120691 341597
rect 127566 341594 127572 341596
rect 120625 341592 127572 341594
rect 120625 341536 120630 341592
rect 120686 341536 127572 341592
rect 120625 341534 127572 341536
rect 120625 341531 120691 341534
rect 127566 341532 127572 341534
rect 127636 341532 127642 341596
rect 135345 341594 135411 341597
rect 164141 341594 164207 341597
rect 135345 341592 164207 341594
rect 135345 341536 135350 341592
rect 135406 341536 164146 341592
rect 164202 341536 164207 341592
rect 135345 341534 164207 341536
rect 135345 341531 135411 341534
rect 164141 341531 164207 341534
rect 90541 341458 90607 341461
rect 322197 341458 322263 341461
rect 326429 341458 326495 341461
rect 328453 341458 328519 341461
rect 90541 341456 322263 341458
rect 90541 341400 90546 341456
rect 90602 341400 322202 341456
rect 322258 341400 322263 341456
rect 90541 341398 322263 341400
rect 90541 341395 90607 341398
rect 322197 341395 322263 341398
rect 325650 341456 326495 341458
rect 325650 341400 326434 341456
rect 326490 341400 326495 341456
rect 325650 341398 326495 341400
rect 90357 341322 90423 341325
rect 325650 341322 325710 341398
rect 326429 341395 326495 341398
rect 327214 341456 328519 341458
rect 327214 341400 328458 341456
rect 328514 341400 328519 341456
rect 327214 341398 328519 341400
rect 90357 341320 325710 341322
rect 90357 341264 90362 341320
rect 90418 341264 325710 341320
rect 90357 341262 325710 341264
rect 90357 341259 90423 341262
rect 3366 341124 3372 341188
rect 3436 341186 3442 341188
rect 327214 341186 327274 341398
rect 328453 341395 328519 341398
rect 330334 341396 330340 341460
rect 330404 341458 330410 341460
rect 330661 341458 330727 341461
rect 330404 341456 330727 341458
rect 330404 341400 330666 341456
rect 330722 341400 330727 341456
rect 330404 341398 330727 341400
rect 330404 341396 330410 341398
rect 330661 341395 330727 341398
rect 3436 341126 327274 341186
rect 3436 341124 3442 341126
rect 127566 340988 127572 341052
rect 127636 341050 127642 341052
rect 580717 341050 580783 341053
rect 127636 341048 580783 341050
rect 127636 340992 580722 341048
rect 580778 340992 580783 341048
rect 127636 340990 580783 340992
rect 127636 340988 127642 340990
rect 580717 340987 580783 340990
rect 110454 340852 110460 340916
rect 110524 340914 110530 340916
rect 580349 340914 580415 340917
rect 110524 340912 580415 340914
rect 110524 340856 580354 340912
rect 580410 340856 580415 340912
rect 110524 340854 580415 340856
rect 110524 340852 110530 340854
rect 580349 340851 580415 340854
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580073 325274 580139 325277
rect 583520 325274 584960 325364
rect 580073 325272 584960 325274
rect 580073 325216 580078 325272
rect 580134 325216 584960 325272
rect 580073 325214 584960 325216
rect 580073 325211 580139 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3233 319290 3299 319293
rect -960 319288 3299 319290
rect -960 319232 3238 319288
rect 3294 319232 3299 319288
rect -960 319230 3299 319232
rect -960 319140 480 319230
rect 3233 319227 3299 319230
rect 583520 312082 584960 312172
rect 567150 312022 584960 312082
rect 328126 311884 328132 311948
rect 328196 311946 328202 311948
rect 567150 311946 567210 312022
rect 328196 311886 567210 311946
rect 583520 311932 584960 312022
rect 328196 311884 328202 311886
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 580901 298754 580967 298757
rect 583520 298754 584960 298844
rect 580901 298752 584960 298754
rect 580901 298696 580906 298752
rect 580962 298696 584960 298752
rect 580901 298694 584960 298696
rect 580901 298691 580967 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 4061 293178 4127 293181
rect -960 293176 4127 293178
rect -960 293120 4066 293176
rect 4122 293120 4127 293176
rect -960 293118 4127 293120
rect -960 293028 480 293118
rect 4061 293115 4127 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272234 584960 272324
rect 567150 272174 584960 272234
rect 329046 271900 329052 271964
rect 329116 271962 329122 271964
rect 567150 271962 567210 272174
rect 583520 272084 584960 272174
rect 329116 271902 567210 271962
rect 329116 271900 329122 271902
rect -960 267202 480 267292
rect 3969 267202 4035 267205
rect -960 267200 4035 267202
rect -960 267144 3974 267200
rect 4030 267144 4035 267200
rect -960 267142 4035 267144
rect -960 267052 480 267142
rect 3969 267139 4035 267142
rect 583520 258906 584960 258996
rect 583342 258846 584960 258906
rect 583342 258770 583402 258846
rect 583520 258770 584960 258846
rect 583342 258756 584960 258770
rect 583342 258710 583586 258756
rect 327942 258028 327948 258092
rect 328012 258028 328018 258092
rect 327950 257954 328010 258028
rect 583526 257954 583586 258710
rect 327950 257894 583586 257954
rect -960 254146 480 254236
rect 3877 254146 3943 254149
rect -960 254144 3943 254146
rect -960 254088 3882 254144
rect 3938 254088 3943 254144
rect -960 254086 3943 254088
rect -960 253996 480 254086
rect 3877 254083 3943 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3785 241090 3851 241093
rect -960 241088 3851 241090
rect -960 241032 3790 241088
rect 3846 241032 3851 241088
rect -960 241030 3851 241032
rect -960 240940 480 241030
rect 3785 241027 3851 241030
rect 580073 232386 580139 232389
rect 583520 232386 584960 232476
rect 580073 232384 584960 232386
rect 580073 232328 580078 232384
rect 580134 232328 584960 232384
rect 580073 232326 584960 232328
rect 580073 232323 580139 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 583520 219058 584960 219148
rect 583342 218998 584960 219058
rect 583342 218922 583402 218998
rect 583520 218922 584960 218998
rect 583342 218908 584960 218922
rect 583342 218862 583586 218908
rect 327758 218044 327764 218108
rect 327828 218106 327834 218108
rect 583526 218106 583586 218862
rect 327828 218046 583586 218106
rect 327828 218044 327834 218046
rect -960 214978 480 215068
rect 3693 214978 3759 214981
rect -960 214976 3759 214978
rect -960 214920 3698 214976
rect 3754 214920 3759 214976
rect -960 214918 3759 214920
rect -960 214828 480 214918
rect 3693 214915 3759 214918
rect 580809 205730 580875 205733
rect 583520 205730 584960 205820
rect 580809 205728 584960 205730
rect 580809 205672 580814 205728
rect 580870 205672 584960 205728
rect 580809 205670 584960 205672
rect 580809 205667 580875 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3601 201922 3667 201925
rect -960 201920 3667 201922
rect -960 201864 3606 201920
rect 3662 201864 3667 201920
rect -960 201862 3667 201864
rect -960 201772 480 201862
rect 3601 201859 3667 201862
rect 580717 192538 580783 192541
rect 583520 192538 584960 192628
rect 580717 192536 584960 192538
rect 580717 192480 580722 192536
rect 580778 192480 584960 192536
rect 580717 192478 584960 192480
rect 580717 192475 580783 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 580625 179210 580691 179213
rect 583520 179210 584960 179300
rect 580625 179208 584960 179210
rect 580625 179152 580630 179208
rect 580686 179152 584960 179208
rect 580625 179150 584960 179152
rect 580625 179147 580691 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580533 165882 580599 165885
rect 583520 165882 584960 165972
rect 580533 165880 584960 165882
rect 580533 165824 580538 165880
rect 580594 165824 584960 165880
rect 580533 165822 584960 165824
rect 580533 165819 580599 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 2773 162890 2839 162893
rect -960 162888 2839 162890
rect -960 162832 2778 162888
rect 2834 162832 2839 162888
rect -960 162830 2839 162832
rect -960 162740 480 162830
rect 2773 162827 2839 162830
rect 580901 152690 580967 152693
rect 583520 152690 584960 152780
rect 580901 152688 584960 152690
rect 580901 152632 580906 152688
rect 580962 152632 584960 152688
rect 580901 152630 584960 152632
rect 580901 152627 580967 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 583520 139362 584960 139452
rect 583342 139302 584960 139362
rect 583342 139226 583402 139302
rect 583520 139226 584960 139302
rect 583342 139212 584960 139226
rect 583342 139166 583586 139212
rect 327574 138076 327580 138140
rect 327644 138138 327650 138140
rect 583526 138138 583586 139166
rect 327644 138078 583586 138138
rect 327644 138076 327650 138078
rect -960 136778 480 136868
rect 3550 136778 3556 136780
rect -960 136718 3556 136778
rect -960 136628 480 136718
rect 3550 136716 3556 136718
rect 3620 136716 3626 136780
rect 580441 126034 580507 126037
rect 583520 126034 584960 126124
rect 580441 126032 584960 126034
rect 580441 125976 580446 126032
rect 580502 125976 584960 126032
rect 580441 125974 584960 125976
rect 580441 125971 580507 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 580349 112842 580415 112845
rect 583520 112842 584960 112932
rect 580349 112840 584960 112842
rect 580349 112784 580354 112840
rect 580410 112784 584960 112840
rect 580349 112782 584960 112784
rect 580349 112779 580415 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 2773 110666 2839 110669
rect -960 110664 2839 110666
rect -960 110608 2778 110664
rect 2834 110608 2839 110664
rect -960 110606 2839 110608
rect -960 110516 480 110606
rect 2773 110603 2839 110606
rect 579981 99514 580047 99517
rect 583520 99514 584960 99604
rect 579981 99512 584960 99514
rect 579981 99456 579986 99512
rect 580042 99456 584960 99512
rect 579981 99454 584960 99456
rect 579981 99451 580047 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 580257 86186 580323 86189
rect 583520 86186 584960 86276
rect 580257 86184 584960 86186
rect 580257 86128 580262 86184
rect 580318 86128 584960 86184
rect 580257 86126 584960 86128
rect 580257 86123 580323 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 579705 72994 579771 72997
rect 583520 72994 584960 73084
rect 579705 72992 584960 72994
rect 579705 72936 579710 72992
rect 579766 72936 584960 72992
rect 579705 72934 584960 72936
rect 579705 72931 579771 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 580206 46276 580212 46340
rect 580276 46338 580282 46340
rect 583520 46338 584960 46428
rect 580276 46278 584960 46338
rect 580276 46276 580282 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 579613 33146 579679 33149
rect 583520 33146 584960 33236
rect 579613 33144 584960 33146
rect 579613 33088 579618 33144
rect 579674 33088 584960 33144
rect 579613 33086 584960 33088
rect 579613 33083 579679 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3141 32466 3207 32469
rect -960 32464 3207 32466
rect -960 32408 3146 32464
rect 3202 32408 3207 32464
rect -960 32406 3207 32408
rect -960 32316 480 32406
rect 3141 32403 3207 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 330334 19410 330340 19412
rect -960 19350 330340 19410
rect -960 19260 480 19350
rect 330334 19348 330340 19350
rect 330404 19348 330410 19412
rect 328637 18594 328703 18597
rect 576853 18594 576919 18597
rect 328637 18592 576919 18594
rect 328637 18536 328642 18592
rect 328698 18536 576858 18592
rect 576914 18536 576919 18592
rect 328637 18534 576919 18536
rect 328637 18531 328703 18534
rect 576853 18531 576919 18534
rect 329925 15874 329991 15877
rect 578601 15874 578667 15877
rect 329925 15872 578667 15874
rect 329925 15816 329930 15872
rect 329986 15816 578606 15872
rect 578662 15816 578667 15872
rect 329925 15814 578667 15816
rect 329925 15811 329991 15814
rect 578601 15811 578667 15814
rect 306557 14514 306623 14517
rect 521653 14514 521719 14517
rect 306557 14512 521719 14514
rect 306557 14456 306562 14512
rect 306618 14456 521658 14512
rect 521714 14456 521719 14512
rect 306557 14454 521719 14456
rect 306557 14451 306623 14454
rect 521653 14451 521719 14454
rect 320265 11658 320331 11661
rect 556153 11658 556219 11661
rect 320265 11656 556219 11658
rect 320265 11600 320270 11656
rect 320326 11600 556158 11656
rect 556214 11600 556219 11656
rect 320265 11598 556219 11600
rect 320265 11595 320331 11598
rect 556153 11595 556219 11598
rect 321553 10298 321619 10301
rect 559281 10298 559347 10301
rect 321553 10296 559347 10298
rect 321553 10240 321558 10296
rect 321614 10240 559286 10296
rect 559342 10240 559347 10296
rect 321553 10238 559347 10240
rect 321553 10235 321619 10238
rect 559281 10235 559347 10238
rect 295333 8938 295399 8941
rect 495893 8938 495959 8941
rect 295333 8936 495959 8938
rect 295333 8880 295338 8936
rect 295394 8880 495898 8936
rect 495954 8880 495959 8936
rect 295333 8878 495959 8880
rect 295333 8875 295399 8878
rect 495893 8875 495959 8878
rect -960 6490 480 6580
rect 580758 6564 580764 6628
rect 580828 6626 580834 6628
rect 583520 6626 584960 6716
rect 580828 6566 584960 6626
rect 580828 6564 580834 6566
rect 3366 6490 3372 6492
rect -960 6430 3372 6490
rect -960 6340 480 6430
rect 3366 6428 3372 6430
rect 3436 6428 3442 6492
rect 583520 6476 584960 6566
rect 13537 6218 13603 6221
rect 96705 6218 96771 6221
rect 13537 6216 96771 6218
rect 13537 6160 13542 6216
rect 13598 6160 96710 6216
rect 96766 6160 96771 6216
rect 13537 6158 96771 6160
rect 13537 6155 13603 6158
rect 96705 6155 96771 6158
rect 236269 6218 236335 6221
rect 352833 6218 352899 6221
rect 236269 6216 352899 6218
rect 236269 6160 236274 6216
rect 236330 6160 352838 6216
rect 352894 6160 352899 6216
rect 236269 6158 352899 6160
rect 236269 6155 236335 6158
rect 352833 6155 352899 6158
rect 65517 4858 65583 4861
rect 118785 4858 118851 4861
rect 65517 4856 118851 4858
rect 65517 4800 65522 4856
rect 65578 4800 118790 4856
rect 118846 4800 118851 4856
rect 65517 4798 118851 4800
rect 65517 4795 65583 4798
rect 118785 4795 118851 4798
rect 219433 4858 219499 4861
rect 310237 4858 310303 4861
rect 219433 4856 310303 4858
rect 219433 4800 219438 4856
rect 219494 4800 310242 4856
rect 310298 4800 310303 4856
rect 219433 4798 310303 4800
rect 219433 4795 219499 4798
rect 310237 4795 310303 4798
rect 311893 4858 311959 4861
rect 537201 4858 537267 4861
rect 311893 4856 537267 4858
rect 311893 4800 311898 4856
rect 311954 4800 537206 4856
rect 537262 4800 537267 4856
rect 311893 4798 537267 4800
rect 311893 4795 311959 4798
rect 537201 4795 537267 4798
rect 5257 3362 5323 3365
rect 94037 3362 94103 3365
rect 5257 3360 94103 3362
rect 5257 3304 5262 3360
rect 5318 3304 94042 3360
rect 94098 3304 94103 3360
rect 5257 3302 94103 3304
rect 5257 3299 5323 3302
rect 94037 3299 94103 3302
rect 109309 3362 109375 3365
rect 136725 3362 136791 3365
rect 109309 3360 136791 3362
rect 109309 3304 109314 3360
rect 109370 3304 136730 3360
rect 136786 3304 136791 3360
rect 109309 3302 136791 3304
rect 109309 3299 109375 3302
rect 136725 3299 136791 3302
rect 406377 3362 406443 3365
rect 583385 3362 583451 3365
rect 406377 3360 583451 3362
rect 406377 3304 406382 3360
rect 406438 3304 583390 3360
rect 583446 3304 583451 3360
rect 406377 3302 583451 3304
rect 406377 3299 406443 3302
rect 583385 3299 583451 3302
<< via3 >>
rect 580212 344660 580276 344724
rect 328132 344524 328196 344588
rect 327948 344388 328012 344452
rect 329052 344252 329116 344316
rect 327764 344116 327828 344180
rect 327580 343980 327644 344044
rect 3556 343844 3620 343908
rect 580764 343708 580828 343772
rect 110460 341532 110524 341596
rect 127572 341532 127636 341596
rect 3372 341124 3436 341188
rect 330340 341396 330404 341460
rect 127572 340988 127636 341052
rect 110460 340852 110524 340916
rect 328132 311884 328196 311948
rect 329052 271900 329116 271964
rect 327948 258028 328012 258092
rect 327764 218044 327828 218108
rect 327580 138076 327644 138140
rect 3556 136716 3620 136780
rect 580212 46276 580276 46340
rect 330340 19348 330404 19412
rect 580764 6564 580828 6628
rect 3372 6428 3436 6492
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 3555 343908 3621 343909
rect 3555 343844 3556 343908
rect 3620 343844 3621 343908
rect 3555 343843 3621 343844
rect 3371 341188 3437 341189
rect 3371 341124 3372 341188
rect 3436 341124 3437 341188
rect 3371 341123 3437 341124
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 3374 6493 3434 341123
rect 3558 136781 3618 343843
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 3555 136780 3621 136781
rect 3555 136716 3556 136780
rect 3620 136716 3621 136780
rect 3555 136715 3621 136716
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 3371 6492 3437 6493
rect 3371 6428 3372 6492
rect 3436 6428 3437 6492
rect 3371 6427 3437 6428
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 344000 92414 344898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 344000 96134 348618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 344000 99854 352338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 344000 103574 356058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 344000 110414 362898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 344000 114134 366618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 344000 117854 370338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 344000 121574 374058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 344000 128414 344898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 344000 132134 348618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 344000 135854 352338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 344000 139574 356058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 344000 146414 362898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 344000 150134 366618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 344000 153854 370338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 344000 157574 374058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 344000 164414 344898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 344000 168134 348618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 344000 171854 352338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 344000 175574 356058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 344000 182414 362898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 344000 186134 366618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 344000 189854 370338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 344000 193574 374058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 344000 200414 344898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 344000 204134 348618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 344000 207854 352338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 344000 211574 356058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 344000 218414 362898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 344000 222134 366618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 344000 225854 370338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 344000 229574 374058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 344000 236414 344898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 344000 240134 348618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 344000 243854 352338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 344000 247574 356058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 344000 254414 362898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 344000 258134 366618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 344000 261854 370338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 344000 265574 374058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 344000 272414 344898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 344000 276134 348618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 344000 279854 352338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 344000 283574 356058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 344000 290414 362898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 344000 294134 366618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 344000 297854 370338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 344000 301574 374058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 344000 308414 344898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 344000 312134 348618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 344000 315854 352338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 344000 319574 356058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 344000 326414 362898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 328131 344588 328197 344589
rect 328131 344524 328132 344588
rect 328196 344524 328197 344588
rect 328131 344523 328197 344524
rect 327947 344452 328013 344453
rect 327947 344388 327948 344452
rect 328012 344388 328013 344452
rect 327947 344387 328013 344388
rect 327763 344180 327829 344181
rect 327763 344116 327764 344180
rect 327828 344116 327829 344180
rect 327763 344115 327829 344116
rect 327579 344044 327645 344045
rect 327579 343980 327580 344044
rect 327644 343980 327645 344044
rect 327579 343979 327645 343980
rect 110459 341596 110525 341597
rect 110459 341532 110460 341596
rect 110524 341532 110525 341596
rect 110459 341531 110525 341532
rect 127571 341596 127637 341597
rect 127571 341532 127572 341596
rect 127636 341532 127637 341596
rect 127571 341531 127637 341532
rect 110462 340917 110522 341531
rect 127574 341053 127634 341531
rect 127571 341052 127637 341053
rect 127571 340988 127572 341052
rect 127636 340988 127637 341052
rect 127571 340987 127637 340988
rect 110459 340916 110525 340917
rect 110459 340852 110460 340916
rect 110524 340852 110525 340916
rect 110459 340851 110525 340852
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 96208 327454 96528 327486
rect 96208 327218 96250 327454
rect 96486 327218 96528 327454
rect 96208 327134 96528 327218
rect 96208 326898 96250 327134
rect 96486 326898 96528 327134
rect 96208 326866 96528 326898
rect 126928 327454 127248 327486
rect 126928 327218 126970 327454
rect 127206 327218 127248 327454
rect 126928 327134 127248 327218
rect 126928 326898 126970 327134
rect 127206 326898 127248 327134
rect 126928 326866 127248 326898
rect 157648 327454 157968 327486
rect 157648 327218 157690 327454
rect 157926 327218 157968 327454
rect 157648 327134 157968 327218
rect 157648 326898 157690 327134
rect 157926 326898 157968 327134
rect 157648 326866 157968 326898
rect 188368 327454 188688 327486
rect 188368 327218 188410 327454
rect 188646 327218 188688 327454
rect 188368 327134 188688 327218
rect 188368 326898 188410 327134
rect 188646 326898 188688 327134
rect 188368 326866 188688 326898
rect 219088 327454 219408 327486
rect 219088 327218 219130 327454
rect 219366 327218 219408 327454
rect 219088 327134 219408 327218
rect 219088 326898 219130 327134
rect 219366 326898 219408 327134
rect 219088 326866 219408 326898
rect 249808 327454 250128 327486
rect 249808 327218 249850 327454
rect 250086 327218 250128 327454
rect 249808 327134 250128 327218
rect 249808 326898 249850 327134
rect 250086 326898 250128 327134
rect 249808 326866 250128 326898
rect 280528 327454 280848 327486
rect 280528 327218 280570 327454
rect 280806 327218 280848 327454
rect 280528 327134 280848 327218
rect 280528 326898 280570 327134
rect 280806 326898 280848 327134
rect 280528 326866 280848 326898
rect 311248 327454 311568 327486
rect 311248 327218 311290 327454
rect 311526 327218 311568 327454
rect 311248 327134 311568 327218
rect 311248 326898 311290 327134
rect 311526 326898 311568 327134
rect 311248 326866 311568 326898
rect 111568 309454 111888 309486
rect 111568 309218 111610 309454
rect 111846 309218 111888 309454
rect 111568 309134 111888 309218
rect 111568 308898 111610 309134
rect 111846 308898 111888 309134
rect 111568 308866 111888 308898
rect 142288 309454 142608 309486
rect 142288 309218 142330 309454
rect 142566 309218 142608 309454
rect 142288 309134 142608 309218
rect 142288 308898 142330 309134
rect 142566 308898 142608 309134
rect 142288 308866 142608 308898
rect 173008 309454 173328 309486
rect 173008 309218 173050 309454
rect 173286 309218 173328 309454
rect 173008 309134 173328 309218
rect 173008 308898 173050 309134
rect 173286 308898 173328 309134
rect 173008 308866 173328 308898
rect 203728 309454 204048 309486
rect 203728 309218 203770 309454
rect 204006 309218 204048 309454
rect 203728 309134 204048 309218
rect 203728 308898 203770 309134
rect 204006 308898 204048 309134
rect 203728 308866 204048 308898
rect 234448 309454 234768 309486
rect 234448 309218 234490 309454
rect 234726 309218 234768 309454
rect 234448 309134 234768 309218
rect 234448 308898 234490 309134
rect 234726 308898 234768 309134
rect 234448 308866 234768 308898
rect 265168 309454 265488 309486
rect 265168 309218 265210 309454
rect 265446 309218 265488 309454
rect 265168 309134 265488 309218
rect 265168 308898 265210 309134
rect 265446 308898 265488 309134
rect 265168 308866 265488 308898
rect 295888 309454 296208 309486
rect 295888 309218 295930 309454
rect 296166 309218 296208 309454
rect 295888 309134 296208 309218
rect 295888 308898 295930 309134
rect 296166 308898 296208 309134
rect 295888 308866 296208 308898
rect 326608 309454 326928 309486
rect 326608 309218 326650 309454
rect 326886 309218 326928 309454
rect 326608 309134 326928 309218
rect 326608 308898 326650 309134
rect 326886 308898 326928 309134
rect 326608 308866 326928 308898
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 96208 291454 96528 291486
rect 96208 291218 96250 291454
rect 96486 291218 96528 291454
rect 96208 291134 96528 291218
rect 96208 290898 96250 291134
rect 96486 290898 96528 291134
rect 96208 290866 96528 290898
rect 126928 291454 127248 291486
rect 126928 291218 126970 291454
rect 127206 291218 127248 291454
rect 126928 291134 127248 291218
rect 126928 290898 126970 291134
rect 127206 290898 127248 291134
rect 126928 290866 127248 290898
rect 157648 291454 157968 291486
rect 157648 291218 157690 291454
rect 157926 291218 157968 291454
rect 157648 291134 157968 291218
rect 157648 290898 157690 291134
rect 157926 290898 157968 291134
rect 157648 290866 157968 290898
rect 188368 291454 188688 291486
rect 188368 291218 188410 291454
rect 188646 291218 188688 291454
rect 188368 291134 188688 291218
rect 188368 290898 188410 291134
rect 188646 290898 188688 291134
rect 188368 290866 188688 290898
rect 219088 291454 219408 291486
rect 219088 291218 219130 291454
rect 219366 291218 219408 291454
rect 219088 291134 219408 291218
rect 219088 290898 219130 291134
rect 219366 290898 219408 291134
rect 219088 290866 219408 290898
rect 249808 291454 250128 291486
rect 249808 291218 249850 291454
rect 250086 291218 250128 291454
rect 249808 291134 250128 291218
rect 249808 290898 249850 291134
rect 250086 290898 250128 291134
rect 249808 290866 250128 290898
rect 280528 291454 280848 291486
rect 280528 291218 280570 291454
rect 280806 291218 280848 291454
rect 280528 291134 280848 291218
rect 280528 290898 280570 291134
rect 280806 290898 280848 291134
rect 280528 290866 280848 290898
rect 311248 291454 311568 291486
rect 311248 291218 311290 291454
rect 311526 291218 311568 291454
rect 311248 291134 311568 291218
rect 311248 290898 311290 291134
rect 311526 290898 311568 291134
rect 311248 290866 311568 290898
rect 111568 273454 111888 273486
rect 111568 273218 111610 273454
rect 111846 273218 111888 273454
rect 111568 273134 111888 273218
rect 111568 272898 111610 273134
rect 111846 272898 111888 273134
rect 111568 272866 111888 272898
rect 142288 273454 142608 273486
rect 142288 273218 142330 273454
rect 142566 273218 142608 273454
rect 142288 273134 142608 273218
rect 142288 272898 142330 273134
rect 142566 272898 142608 273134
rect 142288 272866 142608 272898
rect 173008 273454 173328 273486
rect 173008 273218 173050 273454
rect 173286 273218 173328 273454
rect 173008 273134 173328 273218
rect 173008 272898 173050 273134
rect 173286 272898 173328 273134
rect 173008 272866 173328 272898
rect 203728 273454 204048 273486
rect 203728 273218 203770 273454
rect 204006 273218 204048 273454
rect 203728 273134 204048 273218
rect 203728 272898 203770 273134
rect 204006 272898 204048 273134
rect 203728 272866 204048 272898
rect 234448 273454 234768 273486
rect 234448 273218 234490 273454
rect 234726 273218 234768 273454
rect 234448 273134 234768 273218
rect 234448 272898 234490 273134
rect 234726 272898 234768 273134
rect 234448 272866 234768 272898
rect 265168 273454 265488 273486
rect 265168 273218 265210 273454
rect 265446 273218 265488 273454
rect 265168 273134 265488 273218
rect 265168 272898 265210 273134
rect 265446 272898 265488 273134
rect 265168 272866 265488 272898
rect 295888 273454 296208 273486
rect 295888 273218 295930 273454
rect 296166 273218 296208 273454
rect 295888 273134 296208 273218
rect 295888 272898 295930 273134
rect 296166 272898 296208 273134
rect 295888 272866 296208 272898
rect 326608 273454 326928 273486
rect 326608 273218 326650 273454
rect 326886 273218 326928 273454
rect 326608 273134 326928 273218
rect 326608 272898 326650 273134
rect 326886 272898 326928 273134
rect 326608 272866 326928 272898
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 96208 255454 96528 255486
rect 96208 255218 96250 255454
rect 96486 255218 96528 255454
rect 96208 255134 96528 255218
rect 96208 254898 96250 255134
rect 96486 254898 96528 255134
rect 96208 254866 96528 254898
rect 126928 255454 127248 255486
rect 126928 255218 126970 255454
rect 127206 255218 127248 255454
rect 126928 255134 127248 255218
rect 126928 254898 126970 255134
rect 127206 254898 127248 255134
rect 126928 254866 127248 254898
rect 157648 255454 157968 255486
rect 157648 255218 157690 255454
rect 157926 255218 157968 255454
rect 157648 255134 157968 255218
rect 157648 254898 157690 255134
rect 157926 254898 157968 255134
rect 157648 254866 157968 254898
rect 188368 255454 188688 255486
rect 188368 255218 188410 255454
rect 188646 255218 188688 255454
rect 188368 255134 188688 255218
rect 188368 254898 188410 255134
rect 188646 254898 188688 255134
rect 188368 254866 188688 254898
rect 219088 255454 219408 255486
rect 219088 255218 219130 255454
rect 219366 255218 219408 255454
rect 219088 255134 219408 255218
rect 219088 254898 219130 255134
rect 219366 254898 219408 255134
rect 219088 254866 219408 254898
rect 249808 255454 250128 255486
rect 249808 255218 249850 255454
rect 250086 255218 250128 255454
rect 249808 255134 250128 255218
rect 249808 254898 249850 255134
rect 250086 254898 250128 255134
rect 249808 254866 250128 254898
rect 280528 255454 280848 255486
rect 280528 255218 280570 255454
rect 280806 255218 280848 255454
rect 280528 255134 280848 255218
rect 280528 254898 280570 255134
rect 280806 254898 280848 255134
rect 280528 254866 280848 254898
rect 311248 255454 311568 255486
rect 311248 255218 311290 255454
rect 311526 255218 311568 255454
rect 311248 255134 311568 255218
rect 311248 254898 311290 255134
rect 311526 254898 311568 255134
rect 311248 254866 311568 254898
rect 111568 237454 111888 237486
rect 111568 237218 111610 237454
rect 111846 237218 111888 237454
rect 111568 237134 111888 237218
rect 111568 236898 111610 237134
rect 111846 236898 111888 237134
rect 111568 236866 111888 236898
rect 142288 237454 142608 237486
rect 142288 237218 142330 237454
rect 142566 237218 142608 237454
rect 142288 237134 142608 237218
rect 142288 236898 142330 237134
rect 142566 236898 142608 237134
rect 142288 236866 142608 236898
rect 173008 237454 173328 237486
rect 173008 237218 173050 237454
rect 173286 237218 173328 237454
rect 173008 237134 173328 237218
rect 173008 236898 173050 237134
rect 173286 236898 173328 237134
rect 173008 236866 173328 236898
rect 203728 237454 204048 237486
rect 203728 237218 203770 237454
rect 204006 237218 204048 237454
rect 203728 237134 204048 237218
rect 203728 236898 203770 237134
rect 204006 236898 204048 237134
rect 203728 236866 204048 236898
rect 234448 237454 234768 237486
rect 234448 237218 234490 237454
rect 234726 237218 234768 237454
rect 234448 237134 234768 237218
rect 234448 236898 234490 237134
rect 234726 236898 234768 237134
rect 234448 236866 234768 236898
rect 265168 237454 265488 237486
rect 265168 237218 265210 237454
rect 265446 237218 265488 237454
rect 265168 237134 265488 237218
rect 265168 236898 265210 237134
rect 265446 236898 265488 237134
rect 265168 236866 265488 236898
rect 295888 237454 296208 237486
rect 295888 237218 295930 237454
rect 296166 237218 296208 237454
rect 295888 237134 296208 237218
rect 295888 236898 295930 237134
rect 296166 236898 296208 237134
rect 295888 236866 296208 236898
rect 326608 237454 326928 237486
rect 326608 237218 326650 237454
rect 326886 237218 326928 237454
rect 326608 237134 326928 237218
rect 326608 236898 326650 237134
rect 326886 236898 326928 237134
rect 326608 236866 326928 236898
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 96208 219454 96528 219486
rect 96208 219218 96250 219454
rect 96486 219218 96528 219454
rect 96208 219134 96528 219218
rect 96208 218898 96250 219134
rect 96486 218898 96528 219134
rect 96208 218866 96528 218898
rect 126928 219454 127248 219486
rect 126928 219218 126970 219454
rect 127206 219218 127248 219454
rect 126928 219134 127248 219218
rect 126928 218898 126970 219134
rect 127206 218898 127248 219134
rect 126928 218866 127248 218898
rect 157648 219454 157968 219486
rect 157648 219218 157690 219454
rect 157926 219218 157968 219454
rect 157648 219134 157968 219218
rect 157648 218898 157690 219134
rect 157926 218898 157968 219134
rect 157648 218866 157968 218898
rect 188368 219454 188688 219486
rect 188368 219218 188410 219454
rect 188646 219218 188688 219454
rect 188368 219134 188688 219218
rect 188368 218898 188410 219134
rect 188646 218898 188688 219134
rect 188368 218866 188688 218898
rect 219088 219454 219408 219486
rect 219088 219218 219130 219454
rect 219366 219218 219408 219454
rect 219088 219134 219408 219218
rect 219088 218898 219130 219134
rect 219366 218898 219408 219134
rect 219088 218866 219408 218898
rect 249808 219454 250128 219486
rect 249808 219218 249850 219454
rect 250086 219218 250128 219454
rect 249808 219134 250128 219218
rect 249808 218898 249850 219134
rect 250086 218898 250128 219134
rect 249808 218866 250128 218898
rect 280528 219454 280848 219486
rect 280528 219218 280570 219454
rect 280806 219218 280848 219454
rect 280528 219134 280848 219218
rect 280528 218898 280570 219134
rect 280806 218898 280848 219134
rect 280528 218866 280848 218898
rect 311248 219454 311568 219486
rect 311248 219218 311290 219454
rect 311526 219218 311568 219454
rect 311248 219134 311568 219218
rect 311248 218898 311290 219134
rect 311526 218898 311568 219134
rect 311248 218866 311568 218898
rect 111568 201454 111888 201486
rect 111568 201218 111610 201454
rect 111846 201218 111888 201454
rect 111568 201134 111888 201218
rect 111568 200898 111610 201134
rect 111846 200898 111888 201134
rect 111568 200866 111888 200898
rect 142288 201454 142608 201486
rect 142288 201218 142330 201454
rect 142566 201218 142608 201454
rect 142288 201134 142608 201218
rect 142288 200898 142330 201134
rect 142566 200898 142608 201134
rect 142288 200866 142608 200898
rect 173008 201454 173328 201486
rect 173008 201218 173050 201454
rect 173286 201218 173328 201454
rect 173008 201134 173328 201218
rect 173008 200898 173050 201134
rect 173286 200898 173328 201134
rect 173008 200866 173328 200898
rect 203728 201454 204048 201486
rect 203728 201218 203770 201454
rect 204006 201218 204048 201454
rect 203728 201134 204048 201218
rect 203728 200898 203770 201134
rect 204006 200898 204048 201134
rect 203728 200866 204048 200898
rect 234448 201454 234768 201486
rect 234448 201218 234490 201454
rect 234726 201218 234768 201454
rect 234448 201134 234768 201218
rect 234448 200898 234490 201134
rect 234726 200898 234768 201134
rect 234448 200866 234768 200898
rect 265168 201454 265488 201486
rect 265168 201218 265210 201454
rect 265446 201218 265488 201454
rect 265168 201134 265488 201218
rect 265168 200898 265210 201134
rect 265446 200898 265488 201134
rect 265168 200866 265488 200898
rect 295888 201454 296208 201486
rect 295888 201218 295930 201454
rect 296166 201218 296208 201454
rect 295888 201134 296208 201218
rect 295888 200898 295930 201134
rect 296166 200898 296208 201134
rect 295888 200866 296208 200898
rect 326608 201454 326928 201486
rect 326608 201218 326650 201454
rect 326886 201218 326928 201454
rect 326608 201134 326928 201218
rect 326608 200898 326650 201134
rect 326886 200898 326928 201134
rect 326608 200866 326928 200898
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 96208 183454 96528 183486
rect 96208 183218 96250 183454
rect 96486 183218 96528 183454
rect 96208 183134 96528 183218
rect 96208 182898 96250 183134
rect 96486 182898 96528 183134
rect 96208 182866 96528 182898
rect 126928 183454 127248 183486
rect 126928 183218 126970 183454
rect 127206 183218 127248 183454
rect 126928 183134 127248 183218
rect 126928 182898 126970 183134
rect 127206 182898 127248 183134
rect 126928 182866 127248 182898
rect 157648 183454 157968 183486
rect 157648 183218 157690 183454
rect 157926 183218 157968 183454
rect 157648 183134 157968 183218
rect 157648 182898 157690 183134
rect 157926 182898 157968 183134
rect 157648 182866 157968 182898
rect 188368 183454 188688 183486
rect 188368 183218 188410 183454
rect 188646 183218 188688 183454
rect 188368 183134 188688 183218
rect 188368 182898 188410 183134
rect 188646 182898 188688 183134
rect 188368 182866 188688 182898
rect 219088 183454 219408 183486
rect 219088 183218 219130 183454
rect 219366 183218 219408 183454
rect 219088 183134 219408 183218
rect 219088 182898 219130 183134
rect 219366 182898 219408 183134
rect 219088 182866 219408 182898
rect 249808 183454 250128 183486
rect 249808 183218 249850 183454
rect 250086 183218 250128 183454
rect 249808 183134 250128 183218
rect 249808 182898 249850 183134
rect 250086 182898 250128 183134
rect 249808 182866 250128 182898
rect 280528 183454 280848 183486
rect 280528 183218 280570 183454
rect 280806 183218 280848 183454
rect 280528 183134 280848 183218
rect 280528 182898 280570 183134
rect 280806 182898 280848 183134
rect 280528 182866 280848 182898
rect 311248 183454 311568 183486
rect 311248 183218 311290 183454
rect 311526 183218 311568 183454
rect 311248 183134 311568 183218
rect 311248 182898 311290 183134
rect 311526 182898 311568 183134
rect 311248 182866 311568 182898
rect 111568 165454 111888 165486
rect 111568 165218 111610 165454
rect 111846 165218 111888 165454
rect 111568 165134 111888 165218
rect 111568 164898 111610 165134
rect 111846 164898 111888 165134
rect 111568 164866 111888 164898
rect 142288 165454 142608 165486
rect 142288 165218 142330 165454
rect 142566 165218 142608 165454
rect 142288 165134 142608 165218
rect 142288 164898 142330 165134
rect 142566 164898 142608 165134
rect 142288 164866 142608 164898
rect 173008 165454 173328 165486
rect 173008 165218 173050 165454
rect 173286 165218 173328 165454
rect 173008 165134 173328 165218
rect 173008 164898 173050 165134
rect 173286 164898 173328 165134
rect 173008 164866 173328 164898
rect 203728 165454 204048 165486
rect 203728 165218 203770 165454
rect 204006 165218 204048 165454
rect 203728 165134 204048 165218
rect 203728 164898 203770 165134
rect 204006 164898 204048 165134
rect 203728 164866 204048 164898
rect 234448 165454 234768 165486
rect 234448 165218 234490 165454
rect 234726 165218 234768 165454
rect 234448 165134 234768 165218
rect 234448 164898 234490 165134
rect 234726 164898 234768 165134
rect 234448 164866 234768 164898
rect 265168 165454 265488 165486
rect 265168 165218 265210 165454
rect 265446 165218 265488 165454
rect 265168 165134 265488 165218
rect 265168 164898 265210 165134
rect 265446 164898 265488 165134
rect 265168 164866 265488 164898
rect 295888 165454 296208 165486
rect 295888 165218 295930 165454
rect 296166 165218 296208 165454
rect 295888 165134 296208 165218
rect 295888 164898 295930 165134
rect 296166 164898 296208 165134
rect 295888 164866 296208 164898
rect 326608 165454 326928 165486
rect 326608 165218 326650 165454
rect 326886 165218 326928 165454
rect 326608 165134 326928 165218
rect 326608 164898 326650 165134
rect 326886 164898 326928 165134
rect 326608 164866 326928 164898
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 96208 147454 96528 147486
rect 96208 147218 96250 147454
rect 96486 147218 96528 147454
rect 96208 147134 96528 147218
rect 96208 146898 96250 147134
rect 96486 146898 96528 147134
rect 96208 146866 96528 146898
rect 126928 147454 127248 147486
rect 126928 147218 126970 147454
rect 127206 147218 127248 147454
rect 126928 147134 127248 147218
rect 126928 146898 126970 147134
rect 127206 146898 127248 147134
rect 126928 146866 127248 146898
rect 157648 147454 157968 147486
rect 157648 147218 157690 147454
rect 157926 147218 157968 147454
rect 157648 147134 157968 147218
rect 157648 146898 157690 147134
rect 157926 146898 157968 147134
rect 157648 146866 157968 146898
rect 188368 147454 188688 147486
rect 188368 147218 188410 147454
rect 188646 147218 188688 147454
rect 188368 147134 188688 147218
rect 188368 146898 188410 147134
rect 188646 146898 188688 147134
rect 188368 146866 188688 146898
rect 219088 147454 219408 147486
rect 219088 147218 219130 147454
rect 219366 147218 219408 147454
rect 219088 147134 219408 147218
rect 219088 146898 219130 147134
rect 219366 146898 219408 147134
rect 219088 146866 219408 146898
rect 249808 147454 250128 147486
rect 249808 147218 249850 147454
rect 250086 147218 250128 147454
rect 249808 147134 250128 147218
rect 249808 146898 249850 147134
rect 250086 146898 250128 147134
rect 249808 146866 250128 146898
rect 280528 147454 280848 147486
rect 280528 147218 280570 147454
rect 280806 147218 280848 147454
rect 280528 147134 280848 147218
rect 280528 146898 280570 147134
rect 280806 146898 280848 147134
rect 280528 146866 280848 146898
rect 311248 147454 311568 147486
rect 311248 147218 311290 147454
rect 311526 147218 311568 147454
rect 311248 147134 311568 147218
rect 311248 146898 311290 147134
rect 311526 146898 311568 147134
rect 311248 146866 311568 146898
rect 327582 138141 327642 343979
rect 327766 218109 327826 344115
rect 327950 258093 328010 344387
rect 328134 311949 328194 344523
rect 329051 344316 329117 344317
rect 329051 344252 329052 344316
rect 329116 344252 329117 344316
rect 329051 344251 329117 344252
rect 328131 311948 328197 311949
rect 328131 311884 328132 311948
rect 328196 311884 328197 311948
rect 328131 311883 328197 311884
rect 329054 271965 329114 344251
rect 329514 344000 330134 366618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 344000 333854 370338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 330339 341460 330405 341461
rect 330339 341396 330340 341460
rect 330404 341396 330405 341460
rect 330339 341395 330405 341396
rect 329051 271964 329117 271965
rect 329051 271900 329052 271964
rect 329116 271900 329117 271964
rect 329051 271899 329117 271900
rect 327947 258092 328013 258093
rect 327947 258028 327948 258092
rect 328012 258028 328013 258092
rect 327947 258027 328013 258028
rect 327763 218108 327829 218109
rect 327763 218044 327764 218108
rect 327828 218044 327829 218108
rect 327763 218043 327829 218044
rect 327579 138140 327645 138141
rect 327579 138076 327580 138140
rect 327644 138076 327645 138140
rect 327579 138075 327645 138076
rect 111568 129454 111888 129486
rect 111568 129218 111610 129454
rect 111846 129218 111888 129454
rect 111568 129134 111888 129218
rect 111568 128898 111610 129134
rect 111846 128898 111888 129134
rect 111568 128866 111888 128898
rect 142288 129454 142608 129486
rect 142288 129218 142330 129454
rect 142566 129218 142608 129454
rect 142288 129134 142608 129218
rect 142288 128898 142330 129134
rect 142566 128898 142608 129134
rect 142288 128866 142608 128898
rect 173008 129454 173328 129486
rect 173008 129218 173050 129454
rect 173286 129218 173328 129454
rect 173008 129134 173328 129218
rect 173008 128898 173050 129134
rect 173286 128898 173328 129134
rect 173008 128866 173328 128898
rect 203728 129454 204048 129486
rect 203728 129218 203770 129454
rect 204006 129218 204048 129454
rect 203728 129134 204048 129218
rect 203728 128898 203770 129134
rect 204006 128898 204048 129134
rect 203728 128866 204048 128898
rect 234448 129454 234768 129486
rect 234448 129218 234490 129454
rect 234726 129218 234768 129454
rect 234448 129134 234768 129218
rect 234448 128898 234490 129134
rect 234726 128898 234768 129134
rect 234448 128866 234768 128898
rect 265168 129454 265488 129486
rect 265168 129218 265210 129454
rect 265446 129218 265488 129454
rect 265168 129134 265488 129218
rect 265168 128898 265210 129134
rect 265446 128898 265488 129134
rect 265168 128866 265488 128898
rect 295888 129454 296208 129486
rect 295888 129218 295930 129454
rect 296166 129218 296208 129454
rect 295888 129134 296208 129218
rect 295888 128898 295930 129134
rect 296166 128898 296208 129134
rect 295888 128866 296208 128898
rect 326608 129454 326928 129486
rect 326608 129218 326650 129454
rect 326886 129218 326928 129454
rect 326608 129134 326928 129218
rect 326608 128898 326650 129134
rect 326886 128898 326928 129134
rect 326608 128866 326928 128898
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 96208 111454 96528 111486
rect 96208 111218 96250 111454
rect 96486 111218 96528 111454
rect 96208 111134 96528 111218
rect 96208 110898 96250 111134
rect 96486 110898 96528 111134
rect 96208 110866 96528 110898
rect 126928 111454 127248 111486
rect 126928 111218 126970 111454
rect 127206 111218 127248 111454
rect 126928 111134 127248 111218
rect 126928 110898 126970 111134
rect 127206 110898 127248 111134
rect 126928 110866 127248 110898
rect 157648 111454 157968 111486
rect 157648 111218 157690 111454
rect 157926 111218 157968 111454
rect 157648 111134 157968 111218
rect 157648 110898 157690 111134
rect 157926 110898 157968 111134
rect 157648 110866 157968 110898
rect 188368 111454 188688 111486
rect 188368 111218 188410 111454
rect 188646 111218 188688 111454
rect 188368 111134 188688 111218
rect 188368 110898 188410 111134
rect 188646 110898 188688 111134
rect 188368 110866 188688 110898
rect 219088 111454 219408 111486
rect 219088 111218 219130 111454
rect 219366 111218 219408 111454
rect 219088 111134 219408 111218
rect 219088 110898 219130 111134
rect 219366 110898 219408 111134
rect 219088 110866 219408 110898
rect 249808 111454 250128 111486
rect 249808 111218 249850 111454
rect 250086 111218 250128 111454
rect 249808 111134 250128 111218
rect 249808 110898 249850 111134
rect 250086 110898 250128 111134
rect 249808 110866 250128 110898
rect 280528 111454 280848 111486
rect 280528 111218 280570 111454
rect 280806 111218 280848 111454
rect 280528 111134 280848 111218
rect 280528 110898 280570 111134
rect 280806 110898 280848 111134
rect 280528 110866 280848 110898
rect 311248 111454 311568 111486
rect 311248 111218 311290 111454
rect 311526 111218 311568 111454
rect 311248 111134 311568 111218
rect 311248 110898 311290 111134
rect 311526 110898 311568 111134
rect 311248 110866 311568 110898
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 93454 92414 100000
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 97174 96134 100000
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 100000
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 100000
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 100000
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 79174 114134 100000
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 82894 117854 100000
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 86614 121574 100000
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 93454 128414 100000
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 97174 132134 100000
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 64894 135854 100000
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 100000
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 75454 146414 100000
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 79174 150134 100000
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 82894 153854 100000
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 86614 157574 100000
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 93454 164414 100000
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 97174 168134 100000
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 64894 171854 100000
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 68614 175574 100000
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 75454 182414 100000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 79174 186134 100000
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 82894 189854 100000
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 86614 193574 100000
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 93454 200414 100000
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 97174 204134 100000
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 64894 207854 100000
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 68614 211574 100000
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 100000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 100000
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 82894 225854 100000
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 86614 229574 100000
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 93454 236414 100000
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 97174 240134 100000
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 64894 243854 100000
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 68614 247574 100000
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 75454 254414 100000
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 79174 258134 100000
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 82894 261854 100000
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 86614 265574 100000
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 93454 272414 100000
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 97174 276134 100000
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 64894 279854 100000
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 68614 283574 100000
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 75454 290414 100000
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 79174 294134 100000
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 82894 297854 100000
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 86614 301574 100000
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 93454 308414 100000
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 97174 312134 100000
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 64894 315854 100000
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 68614 319574 100000
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 75454 326414 100000
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 79174 330134 100000
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 330342 19413 330402 341395
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 333234 82894 333854 100000
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 330339 19412 330405 19413
rect 330339 19348 330340 19412
rect 330404 19348 330405 19412
rect 330339 19347 330405 19348
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 580211 344724 580277 344725
rect 580211 344660 580212 344724
rect 580276 344660 580277 344724
rect 580211 344659 580277 344660
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 580214 46341 580274 344659
rect 580763 343772 580829 343773
rect 580763 343708 580764 343772
rect 580828 343708 580829 343772
rect 580763 343707 580829 343708
rect 580211 46340 580277 46341
rect 580211 46276 580212 46340
rect 580276 46276 580277 46340
rect 580211 46275 580277 46276
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 580766 6629 580826 343707
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 580763 6628 580829 6629
rect 580763 6564 580764 6628
rect 580828 6564 580829 6628
rect 580763 6563 580829 6564
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 96250 327218 96486 327454
rect 96250 326898 96486 327134
rect 126970 327218 127206 327454
rect 126970 326898 127206 327134
rect 157690 327218 157926 327454
rect 157690 326898 157926 327134
rect 188410 327218 188646 327454
rect 188410 326898 188646 327134
rect 219130 327218 219366 327454
rect 219130 326898 219366 327134
rect 249850 327218 250086 327454
rect 249850 326898 250086 327134
rect 280570 327218 280806 327454
rect 280570 326898 280806 327134
rect 311290 327218 311526 327454
rect 311290 326898 311526 327134
rect 111610 309218 111846 309454
rect 111610 308898 111846 309134
rect 142330 309218 142566 309454
rect 142330 308898 142566 309134
rect 173050 309218 173286 309454
rect 173050 308898 173286 309134
rect 203770 309218 204006 309454
rect 203770 308898 204006 309134
rect 234490 309218 234726 309454
rect 234490 308898 234726 309134
rect 265210 309218 265446 309454
rect 265210 308898 265446 309134
rect 295930 309218 296166 309454
rect 295930 308898 296166 309134
rect 326650 309218 326886 309454
rect 326650 308898 326886 309134
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 96250 291218 96486 291454
rect 96250 290898 96486 291134
rect 126970 291218 127206 291454
rect 126970 290898 127206 291134
rect 157690 291218 157926 291454
rect 157690 290898 157926 291134
rect 188410 291218 188646 291454
rect 188410 290898 188646 291134
rect 219130 291218 219366 291454
rect 219130 290898 219366 291134
rect 249850 291218 250086 291454
rect 249850 290898 250086 291134
rect 280570 291218 280806 291454
rect 280570 290898 280806 291134
rect 311290 291218 311526 291454
rect 311290 290898 311526 291134
rect 111610 273218 111846 273454
rect 111610 272898 111846 273134
rect 142330 273218 142566 273454
rect 142330 272898 142566 273134
rect 173050 273218 173286 273454
rect 173050 272898 173286 273134
rect 203770 273218 204006 273454
rect 203770 272898 204006 273134
rect 234490 273218 234726 273454
rect 234490 272898 234726 273134
rect 265210 273218 265446 273454
rect 265210 272898 265446 273134
rect 295930 273218 296166 273454
rect 295930 272898 296166 273134
rect 326650 273218 326886 273454
rect 326650 272898 326886 273134
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 96250 255218 96486 255454
rect 96250 254898 96486 255134
rect 126970 255218 127206 255454
rect 126970 254898 127206 255134
rect 157690 255218 157926 255454
rect 157690 254898 157926 255134
rect 188410 255218 188646 255454
rect 188410 254898 188646 255134
rect 219130 255218 219366 255454
rect 219130 254898 219366 255134
rect 249850 255218 250086 255454
rect 249850 254898 250086 255134
rect 280570 255218 280806 255454
rect 280570 254898 280806 255134
rect 311290 255218 311526 255454
rect 311290 254898 311526 255134
rect 111610 237218 111846 237454
rect 111610 236898 111846 237134
rect 142330 237218 142566 237454
rect 142330 236898 142566 237134
rect 173050 237218 173286 237454
rect 173050 236898 173286 237134
rect 203770 237218 204006 237454
rect 203770 236898 204006 237134
rect 234490 237218 234726 237454
rect 234490 236898 234726 237134
rect 265210 237218 265446 237454
rect 265210 236898 265446 237134
rect 295930 237218 296166 237454
rect 295930 236898 296166 237134
rect 326650 237218 326886 237454
rect 326650 236898 326886 237134
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 96250 219218 96486 219454
rect 96250 218898 96486 219134
rect 126970 219218 127206 219454
rect 126970 218898 127206 219134
rect 157690 219218 157926 219454
rect 157690 218898 157926 219134
rect 188410 219218 188646 219454
rect 188410 218898 188646 219134
rect 219130 219218 219366 219454
rect 219130 218898 219366 219134
rect 249850 219218 250086 219454
rect 249850 218898 250086 219134
rect 280570 219218 280806 219454
rect 280570 218898 280806 219134
rect 311290 219218 311526 219454
rect 311290 218898 311526 219134
rect 111610 201218 111846 201454
rect 111610 200898 111846 201134
rect 142330 201218 142566 201454
rect 142330 200898 142566 201134
rect 173050 201218 173286 201454
rect 173050 200898 173286 201134
rect 203770 201218 204006 201454
rect 203770 200898 204006 201134
rect 234490 201218 234726 201454
rect 234490 200898 234726 201134
rect 265210 201218 265446 201454
rect 265210 200898 265446 201134
rect 295930 201218 296166 201454
rect 295930 200898 296166 201134
rect 326650 201218 326886 201454
rect 326650 200898 326886 201134
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 96250 183218 96486 183454
rect 96250 182898 96486 183134
rect 126970 183218 127206 183454
rect 126970 182898 127206 183134
rect 157690 183218 157926 183454
rect 157690 182898 157926 183134
rect 188410 183218 188646 183454
rect 188410 182898 188646 183134
rect 219130 183218 219366 183454
rect 219130 182898 219366 183134
rect 249850 183218 250086 183454
rect 249850 182898 250086 183134
rect 280570 183218 280806 183454
rect 280570 182898 280806 183134
rect 311290 183218 311526 183454
rect 311290 182898 311526 183134
rect 111610 165218 111846 165454
rect 111610 164898 111846 165134
rect 142330 165218 142566 165454
rect 142330 164898 142566 165134
rect 173050 165218 173286 165454
rect 173050 164898 173286 165134
rect 203770 165218 204006 165454
rect 203770 164898 204006 165134
rect 234490 165218 234726 165454
rect 234490 164898 234726 165134
rect 265210 165218 265446 165454
rect 265210 164898 265446 165134
rect 295930 165218 296166 165454
rect 295930 164898 296166 165134
rect 326650 165218 326886 165454
rect 326650 164898 326886 165134
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 96250 147218 96486 147454
rect 96250 146898 96486 147134
rect 126970 147218 127206 147454
rect 126970 146898 127206 147134
rect 157690 147218 157926 147454
rect 157690 146898 157926 147134
rect 188410 147218 188646 147454
rect 188410 146898 188646 147134
rect 219130 147218 219366 147454
rect 219130 146898 219366 147134
rect 249850 147218 250086 147454
rect 249850 146898 250086 147134
rect 280570 147218 280806 147454
rect 280570 146898 280806 147134
rect 311290 147218 311526 147454
rect 311290 146898 311526 147134
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 111610 129218 111846 129454
rect 111610 128898 111846 129134
rect 142330 129218 142566 129454
rect 142330 128898 142566 129134
rect 173050 129218 173286 129454
rect 173050 128898 173286 129134
rect 203770 129218 204006 129454
rect 203770 128898 204006 129134
rect 234490 129218 234726 129454
rect 234490 128898 234726 129134
rect 265210 129218 265446 129454
rect 265210 128898 265446 129134
rect 295930 129218 296166 129454
rect 295930 128898 296166 129134
rect 326650 129218 326886 129454
rect 326650 128898 326886 129134
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 96250 111218 96486 111454
rect 96250 110898 96486 111134
rect 126970 111218 127206 111454
rect 126970 110898 127206 111134
rect 157690 111218 157926 111454
rect 157690 110898 157926 111134
rect 188410 111218 188646 111454
rect 188410 110898 188646 111134
rect 219130 111218 219366 111454
rect 219130 110898 219366 111134
rect 249850 111218 250086 111454
rect 249850 110898 250086 111134
rect 280570 111218 280806 111454
rect 280570 110898 280806 111134
rect 311290 111218 311526 111454
rect 311290 110898 311526 111134
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 96250 327454
rect 96486 327218 126970 327454
rect 127206 327218 157690 327454
rect 157926 327218 188410 327454
rect 188646 327218 219130 327454
rect 219366 327218 249850 327454
rect 250086 327218 280570 327454
rect 280806 327218 311290 327454
rect 311526 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 96250 327134
rect 96486 326898 126970 327134
rect 127206 326898 157690 327134
rect 157926 326898 188410 327134
rect 188646 326898 219130 327134
rect 219366 326898 249850 327134
rect 250086 326898 280570 327134
rect 280806 326898 311290 327134
rect 311526 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 111610 309454
rect 111846 309218 142330 309454
rect 142566 309218 173050 309454
rect 173286 309218 203770 309454
rect 204006 309218 234490 309454
rect 234726 309218 265210 309454
rect 265446 309218 295930 309454
rect 296166 309218 326650 309454
rect 326886 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 111610 309134
rect 111846 308898 142330 309134
rect 142566 308898 173050 309134
rect 173286 308898 203770 309134
rect 204006 308898 234490 309134
rect 234726 308898 265210 309134
rect 265446 308898 295930 309134
rect 296166 308898 326650 309134
rect 326886 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 96250 291454
rect 96486 291218 126970 291454
rect 127206 291218 157690 291454
rect 157926 291218 188410 291454
rect 188646 291218 219130 291454
rect 219366 291218 249850 291454
rect 250086 291218 280570 291454
rect 280806 291218 311290 291454
rect 311526 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 96250 291134
rect 96486 290898 126970 291134
rect 127206 290898 157690 291134
rect 157926 290898 188410 291134
rect 188646 290898 219130 291134
rect 219366 290898 249850 291134
rect 250086 290898 280570 291134
rect 280806 290898 311290 291134
rect 311526 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 111610 273454
rect 111846 273218 142330 273454
rect 142566 273218 173050 273454
rect 173286 273218 203770 273454
rect 204006 273218 234490 273454
rect 234726 273218 265210 273454
rect 265446 273218 295930 273454
rect 296166 273218 326650 273454
rect 326886 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 111610 273134
rect 111846 272898 142330 273134
rect 142566 272898 173050 273134
rect 173286 272898 203770 273134
rect 204006 272898 234490 273134
rect 234726 272898 265210 273134
rect 265446 272898 295930 273134
rect 296166 272898 326650 273134
rect 326886 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 96250 255454
rect 96486 255218 126970 255454
rect 127206 255218 157690 255454
rect 157926 255218 188410 255454
rect 188646 255218 219130 255454
rect 219366 255218 249850 255454
rect 250086 255218 280570 255454
rect 280806 255218 311290 255454
rect 311526 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 96250 255134
rect 96486 254898 126970 255134
rect 127206 254898 157690 255134
rect 157926 254898 188410 255134
rect 188646 254898 219130 255134
rect 219366 254898 249850 255134
rect 250086 254898 280570 255134
rect 280806 254898 311290 255134
rect 311526 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 111610 237454
rect 111846 237218 142330 237454
rect 142566 237218 173050 237454
rect 173286 237218 203770 237454
rect 204006 237218 234490 237454
rect 234726 237218 265210 237454
rect 265446 237218 295930 237454
rect 296166 237218 326650 237454
rect 326886 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 111610 237134
rect 111846 236898 142330 237134
rect 142566 236898 173050 237134
rect 173286 236898 203770 237134
rect 204006 236898 234490 237134
rect 234726 236898 265210 237134
rect 265446 236898 295930 237134
rect 296166 236898 326650 237134
rect 326886 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 96250 219454
rect 96486 219218 126970 219454
rect 127206 219218 157690 219454
rect 157926 219218 188410 219454
rect 188646 219218 219130 219454
rect 219366 219218 249850 219454
rect 250086 219218 280570 219454
rect 280806 219218 311290 219454
rect 311526 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 96250 219134
rect 96486 218898 126970 219134
rect 127206 218898 157690 219134
rect 157926 218898 188410 219134
rect 188646 218898 219130 219134
rect 219366 218898 249850 219134
rect 250086 218898 280570 219134
rect 280806 218898 311290 219134
rect 311526 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 111610 201454
rect 111846 201218 142330 201454
rect 142566 201218 173050 201454
rect 173286 201218 203770 201454
rect 204006 201218 234490 201454
rect 234726 201218 265210 201454
rect 265446 201218 295930 201454
rect 296166 201218 326650 201454
rect 326886 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 111610 201134
rect 111846 200898 142330 201134
rect 142566 200898 173050 201134
rect 173286 200898 203770 201134
rect 204006 200898 234490 201134
rect 234726 200898 265210 201134
rect 265446 200898 295930 201134
rect 296166 200898 326650 201134
rect 326886 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 96250 183454
rect 96486 183218 126970 183454
rect 127206 183218 157690 183454
rect 157926 183218 188410 183454
rect 188646 183218 219130 183454
rect 219366 183218 249850 183454
rect 250086 183218 280570 183454
rect 280806 183218 311290 183454
rect 311526 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 96250 183134
rect 96486 182898 126970 183134
rect 127206 182898 157690 183134
rect 157926 182898 188410 183134
rect 188646 182898 219130 183134
rect 219366 182898 249850 183134
rect 250086 182898 280570 183134
rect 280806 182898 311290 183134
rect 311526 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 111610 165454
rect 111846 165218 142330 165454
rect 142566 165218 173050 165454
rect 173286 165218 203770 165454
rect 204006 165218 234490 165454
rect 234726 165218 265210 165454
rect 265446 165218 295930 165454
rect 296166 165218 326650 165454
rect 326886 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 111610 165134
rect 111846 164898 142330 165134
rect 142566 164898 173050 165134
rect 173286 164898 203770 165134
rect 204006 164898 234490 165134
rect 234726 164898 265210 165134
rect 265446 164898 295930 165134
rect 296166 164898 326650 165134
rect 326886 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 96250 147454
rect 96486 147218 126970 147454
rect 127206 147218 157690 147454
rect 157926 147218 188410 147454
rect 188646 147218 219130 147454
rect 219366 147218 249850 147454
rect 250086 147218 280570 147454
rect 280806 147218 311290 147454
rect 311526 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 96250 147134
rect 96486 146898 126970 147134
rect 127206 146898 157690 147134
rect 157926 146898 188410 147134
rect 188646 146898 219130 147134
rect 219366 146898 249850 147134
rect 250086 146898 280570 147134
rect 280806 146898 311290 147134
rect 311526 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 111610 129454
rect 111846 129218 142330 129454
rect 142566 129218 173050 129454
rect 173286 129218 203770 129454
rect 204006 129218 234490 129454
rect 234726 129218 265210 129454
rect 265446 129218 295930 129454
rect 296166 129218 326650 129454
rect 326886 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 111610 129134
rect 111846 128898 142330 129134
rect 142566 128898 173050 129134
rect 173286 128898 203770 129134
rect 204006 128898 234490 129134
rect 234726 128898 265210 129134
rect 265446 128898 295930 129134
rect 296166 128898 326650 129134
rect 326886 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 96250 111454
rect 96486 111218 126970 111454
rect 127206 111218 157690 111454
rect 157926 111218 188410 111454
rect 188646 111218 219130 111454
rect 219366 111218 249850 111454
rect 250086 111218 280570 111454
rect 280806 111218 311290 111454
rect 311526 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 96250 111134
rect 96486 110898 126970 111134
rect 127206 110898 157690 111134
rect 157926 110898 188410 111134
rect 188646 110898 219130 111134
rect 219366 110898 249850 111134
rect 250086 110898 280570 111134
rect 280806 110898 311290 111134
rect 311526 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_proj_example  mprj
timestamp 0
transform 1 0 92000 0 1 102000
box 202 0 239738 240000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 100000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 100000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 100000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 100000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 100000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 100000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 100000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 344000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 344000 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 344000 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 344000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 344000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 344000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 344000 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 100000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 100000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 100000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 100000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 100000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 100000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 100000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 344000 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 344000 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 344000 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 344000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 344000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 344000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 344000 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 100000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 100000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 100000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 100000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 100000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 100000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 100000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 344000 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 344000 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 344000 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 344000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 344000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 344000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 344000 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 100000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 100000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 100000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 100000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 100000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 100000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 344000 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 344000 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 344000 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 344000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 344000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 344000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 100000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 100000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 100000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 100000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 100000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 100000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 100000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 344000 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 344000 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 344000 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 344000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 344000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 344000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 344000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 100000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 100000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 100000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 100000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 100000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 100000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 100000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 344000 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 344000 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 344000 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 344000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 344000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 344000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 344000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 100000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 100000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 100000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 100000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 100000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 100000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 100000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 344000 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 344000 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 344000 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 344000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 344000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 344000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 344000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 100000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 100000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 100000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 100000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 100000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 100000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 100000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 344000 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 344000 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 344000 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 344000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 344000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 344000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 344000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
